MACRO MAS0
   SIZE 0.01 BY 0.01 ;
END MAS0

MACRO MAS1
   SIZE 0.02 BY 0.16 ;
END MAS1

MACRO MAS2
   SIZE 0.02 BY 0.16 ;
END MAS2

MACRO MAS3
   SIZE 0.02 BY 0.16 ;
END MAS3

MACRO MAS4
   SIZE 0.04 BY 0.16 ;
END MAS4

MACRO MAS5
   SIZE 0.04 BY 0.16 ;
END MAS5

MACRO MAS6
   SIZE 0.04 BY 0.16 ;
END MAS6

MACRO MAS7
   SIZE 0.04 BY 0.16 ;
END MAS7

MACRO MAS8
   SIZE 0.04 BY 0.16 ;
END MAS8

MACRO MAS9
   SIZE 0.04 BY 0.16 ;
END MAS9

MACRO MAS10
   SIZE 0.04 BY 0.16 ;
END MAS10

MACRO MAS11
   SIZE 0.04 BY 0.16 ;
END MAS11

MACRO MAS12
   SIZE 0.04 BY 0.16 ;
END MAS12

MACRO MAS13
   SIZE 0.06 BY 0.16 ;
END MAS13

MACRO MAS14
   SIZE 0.06 BY 0.16 ;
END MAS14

MACRO MAS15
   SIZE 0.06 BY 0.16 ;
END MAS15

MACRO MAS16
   SIZE 0.06 BY 0.16 ;
END MAS16

MACRO MAS17
   SIZE 0.06 BY 0.16 ;
END MAS17

MACRO MAS18
   SIZE 0.06 BY 0.16 ;
END MAS18

MACRO MAS19
   SIZE 0.06 BY 0.16 ;
END MAS19

MACRO MAS20
   SIZE 0.06 BY 0.16 ;
END MAS20

MACRO MAS21
   SIZE 0.06 BY 0.16 ;
END MAS21

MACRO MAS22
   SIZE 0.06 BY 0.16 ;
END MAS22

MACRO MAS23
   SIZE 0.06 BY 0.16 ;
END MAS23

MACRO MAS24
   SIZE 0.06 BY 0.16 ;
END MAS24

MACRO MAS25
   SIZE 0.06 BY 0.16 ;
END MAS25

MACRO MAS26
   SIZE 0.06 BY 0.16 ;
END MAS26

MACRO MAS27
   SIZE 0.06 BY 0.16 ;
END MAS27

MACRO MAS28
   SIZE 0.06 BY 0.16 ;
END MAS28

MACRO MAS29
   SIZE 0.06 BY 0.16 ;
END MAS29

MACRO MAS30
   SIZE 0.06 BY 0.16 ;
END MAS30

MACRO MAS31
   SIZE 0.06 BY 0.16 ;
END MAS31

MACRO MAS32
   SIZE 0.06 BY 0.16 ;
END MAS32

MACRO MAS33
   SIZE 0.06 BY 0.16 ;
END MAS33

MACRO MAS34
   SIZE 0.06 BY 0.16 ;
END MAS34

MACRO MAS35
   SIZE 0.06 BY 0.16 ;
END MAS35

MACRO MAS36
   SIZE 0.06 BY 0.16 ;
END MAS36

MACRO MAS37
   SIZE 0.06 BY 0.16 ;
END MAS37

MACRO MAS38
   SIZE 0.06 BY 0.16 ;
END MAS38

MACRO MAS39
   SIZE 0.06 BY 0.16 ;
END MAS39

MACRO MAS40
   SIZE 0.06 BY 0.16 ;
END MAS40

MACRO MAS41
   SIZE 0.06 BY 0.16 ;
END MAS41

MACRO MAS42
   SIZE 0.06 BY 0.16 ;
END MAS42

MACRO MAS43
   SIZE 0.06 BY 0.16 ;
END MAS43

MACRO MAS44
   SIZE 0.06 BY 0.16 ;
END MAS44

MACRO MAS45
   SIZE 0.08 BY 0.16 ;
END MAS45

MACRO MAS46
   SIZE 0.08 BY 0.16 ;
END MAS46

MACRO MAS47
   SIZE 0.08 BY 0.16 ;
END MAS47

MACRO MAS48
   SIZE 0.08 BY 0.16 ;
END MAS48

MACRO MAS49
   SIZE 0.08 BY 0.16 ;
END MAS49

MACRO MAS50
   SIZE 0.08 BY 0.16 ;
END MAS50

MACRO MAS51
   SIZE 0.08 BY 0.16 ;
END MAS51

MACRO MAS52
   SIZE 0.08 BY 0.16 ;
END MAS52

MACRO MAS53
   SIZE 0.08 BY 0.16 ;
END MAS53

MACRO MAS54
   SIZE 0.08 BY 0.16 ;
END MAS54

MACRO MAS55
   SIZE 0.08 BY 0.16 ;
END MAS55

MACRO MAS56
   SIZE 0.08 BY 0.16 ;
END MAS56

MACRO MAS57
   SIZE 0.08 BY 0.16 ;
END MAS57

MACRO MAS58
   SIZE 0.08 BY 0.16 ;
END MAS58

MACRO MAS59
   SIZE 0.08 BY 0.16 ;
END MAS59

MACRO MAS60
   SIZE 0.08 BY 0.16 ;
END MAS60

MACRO MAS61
   SIZE 0.08 BY 0.16 ;
END MAS61

MACRO MAS62
   SIZE 0.08 BY 0.16 ;
END MAS62

MACRO MAS63
   SIZE 0.08 BY 0.16 ;
END MAS63

MACRO MAS64
   SIZE 0.08 BY 0.16 ;
END MAS64

MACRO MAS65
   SIZE 0.08 BY 0.16 ;
END MAS65

MACRO MAS66
   SIZE 0.08 BY 0.16 ;
END MAS66

MACRO MAS67
   SIZE 0.08 BY 0.16 ;
END MAS67

MACRO MAS68
   SIZE 0.08 BY 0.16 ;
END MAS68

MACRO MAS69
   SIZE 0.08 BY 0.16 ;
END MAS69

MACRO MAS70
   SIZE 0.08 BY 0.16 ;
END MAS70

MACRO MAS71
   SIZE 0.08 BY 0.16 ;
END MAS71

MACRO MAS72
   SIZE 0.08 BY 0.16 ;
END MAS72

MACRO MAS73
   SIZE 0.08 BY 0.16 ;
END MAS73

MACRO MAS74
   SIZE 0.08 BY 0.16 ;
END MAS74

MACRO MAS75
   SIZE 0.08 BY 0.16 ;
END MAS75

MACRO MAS76
   SIZE 0.08 BY 0.16 ;
END MAS76

MACRO MAS77
   SIZE 0.08 BY 0.16 ;
END MAS77

MACRO MAS78
   SIZE 0.08 BY 0.16 ;
END MAS78

MACRO MAS79
   SIZE 0.08 BY 0.16 ;
END MAS79

MACRO MAS80
   SIZE 0.08 BY 0.16 ;
END MAS80

MACRO MAS81
   SIZE 0.08 BY 0.16 ;
END MAS81

MACRO MAS82
   SIZE 0.08 BY 0.16 ;
END MAS82

MACRO MAS83
   SIZE 0.08 BY 0.16 ;
END MAS83

MACRO MAS84
   SIZE 0.08 BY 0.16 ;
END MAS84

MACRO MAS85
   SIZE 0.08 BY 0.16 ;
END MAS85

MACRO MAS86
   SIZE 0.08 BY 0.16 ;
END MAS86

MACRO MAS87
   SIZE 0.08 BY 0.16 ;
END MAS87

MACRO MAS88
   SIZE 0.08 BY 0.16 ;
END MAS88

MACRO MAS89
   SIZE 0.08 BY 0.16 ;
END MAS89

MACRO MAS90
   SIZE 0.08 BY 0.16 ;
END MAS90

MACRO MAS91
   SIZE 0.08 BY 0.16 ;
END MAS91

MACRO MAS92
   SIZE 0.08 BY 0.16 ;
END MAS92

MACRO MAS93
   SIZE 0.08 BY 0.16 ;
END MAS93

MACRO MAS94
   SIZE 0.08 BY 0.16 ;
END MAS94

MACRO MAS95
   SIZE 0.08 BY 0.16 ;
END MAS95

MACRO MAS96
   SIZE 0.08 BY 0.16 ;
END MAS96

MACRO MAS97
   SIZE 0.08 BY 0.16 ;
END MAS97

MACRO MAS98
   SIZE 0.08 BY 0.16 ;
END MAS98

MACRO MAS99
   SIZE 0.08 BY 0.16 ;
END MAS99

MACRO MAS100
   SIZE 0.08 BY 0.16 ;
END MAS100

MACRO MAS101
   SIZE 0.08 BY 0.16 ;
END MAS101

MACRO MAS102
   SIZE 0.08 BY 0.16 ;
END MAS102

MACRO MAS103
   SIZE 0.08 BY 0.16 ;
END MAS103

MACRO MAS104
   SIZE 0.08 BY 0.16 ;
END MAS104

MACRO MAS105
   SIZE 0.08 BY 0.16 ;
END MAS105

MACRO MAS106
   SIZE 0.08 BY 0.16 ;
END MAS106

MACRO MAS107
   SIZE 0.08 BY 0.16 ;
END MAS107

MACRO MAS108
   SIZE 0.08 BY 0.16 ;
END MAS108

MACRO MAS109
   SIZE 0.08 BY 0.16 ;
END MAS109

MACRO MAS110
   SIZE 0.08 BY 0.16 ;
END MAS110

MACRO MAS111
   SIZE 0.08 BY 0.16 ;
END MAS111

MACRO MAS112
   SIZE 0.08 BY 0.16 ;
END MAS112

MACRO MAS113
   SIZE 0.08 BY 0.16 ;
END MAS113

MACRO MAS114
   SIZE 0.08 BY 0.16 ;
END MAS114

MACRO MAS115
   SIZE 0.08 BY 0.16 ;
END MAS115

MACRO MAS116
   SIZE 0.08 BY 0.16 ;
END MAS116

MACRO MAS117
   SIZE 0.08 BY 0.16 ;
END MAS117

MACRO MAS118
   SIZE 0.08 BY 0.16 ;
END MAS118

MACRO MAS119
   SIZE 0.08 BY 0.16 ;
END MAS119

MACRO MAS120
   SIZE 0.08 BY 0.16 ;
END MAS120

MACRO MAS121
   SIZE 0.08 BY 0.16 ;
END MAS121

MACRO MAS122
   SIZE 0.08 BY 0.16 ;
END MAS122

MACRO MAS123
   SIZE 0.08 BY 0.16 ;
END MAS123

MACRO MAS124
   SIZE 0.08 BY 0.16 ;
END MAS124

MACRO MAS125
   SIZE 0.08 BY 0.16 ;
END MAS125

MACRO MAS126
   SIZE 0.08 BY 0.16 ;
END MAS126

MACRO MAS127
   SIZE 0.08 BY 0.16 ;
END MAS127

MACRO MAS128
   SIZE 0.08 BY 0.16 ;
END MAS128

MACRO MAS129
   SIZE 0.08 BY 0.16 ;
END MAS129

MACRO MAS130
   SIZE 0.08 BY 0.16 ;
END MAS130

MACRO MAS131
   SIZE 0.08 BY 0.16 ;
END MAS131

MACRO MAS132
   SIZE 0.08 BY 0.16 ;
END MAS132

MACRO MAS133
   SIZE 0.08 BY 0.16 ;
END MAS133

MACRO MAS134
   SIZE 0.08 BY 0.16 ;
END MAS134

MACRO MAS135
   SIZE 0.08 BY 0.16 ;
END MAS135

MACRO MAS136
   SIZE 0.08 BY 0.16 ;
END MAS136

MACRO MAS137
   SIZE 0.08 BY 0.16 ;
END MAS137

MACRO MAS138
   SIZE 0.08 BY 0.16 ;
END MAS138

MACRO MAS139
   SIZE 0.08 BY 0.16 ;
END MAS139

MACRO MAS140
   SIZE 0.08 BY 0.16 ;
END MAS140

MACRO MAS141
   SIZE 0.08 BY 0.16 ;
END MAS141

MACRO MAS142
   SIZE 0.08 BY 0.16 ;
END MAS142

MACRO MAS143
   SIZE 0.08 BY 0.16 ;
END MAS143

MACRO MAS144
   SIZE 0.08 BY 0.16 ;
END MAS144

MACRO MAS145
   SIZE 0.08 BY 0.16 ;
END MAS145

MACRO MAS146
   SIZE 0.08 BY 0.16 ;
END MAS146

MACRO MAS147
   SIZE 0.08 BY 0.16 ;
END MAS147

MACRO MAS148
   SIZE 0.08 BY 0.16 ;
END MAS148

MACRO MAS149
   SIZE 0.08 BY 0.16 ;
END MAS149

MACRO MAS150
   SIZE 0.08 BY 0.16 ;
END MAS150

MACRO MAS151
   SIZE 0.08 BY 0.16 ;
END MAS151

MACRO MAS152
   SIZE 0.08 BY 0.16 ;
END MAS152

MACRO MAS153
   SIZE 0.08 BY 0.16 ;
END MAS153

MACRO MAS154
   SIZE 0.08 BY 0.16 ;
END MAS154

MACRO MAS155
   SIZE 0.08 BY 0.16 ;
END MAS155

MACRO MAS156
   SIZE 0.08 BY 0.16 ;
END MAS156

MACRO MAS157
   SIZE 0.08 BY 0.16 ;
END MAS157

MACRO MAS158
   SIZE 0.08 BY 0.16 ;
END MAS158

MACRO MAS159
   SIZE 0.08 BY 0.16 ;
END MAS159

MACRO MAS160
   SIZE 0.08 BY 0.16 ;
END MAS160

MACRO MAS161
   SIZE 0.08 BY 0.16 ;
END MAS161

MACRO MAS162
   SIZE 0.08 BY 0.16 ;
END MAS162

MACRO MAS163
   SIZE 0.08 BY 0.16 ;
END MAS163

MACRO MAS164
   SIZE 0.08 BY 0.16 ;
END MAS164

MACRO MAS165
   SIZE 0.08 BY 0.16 ;
END MAS165

MACRO MAS166
   SIZE 0.08 BY 0.16 ;
END MAS166

MACRO MAS167
   SIZE 0.08 BY 0.16 ;
END MAS167

MACRO MAS168
   SIZE 0.08 BY 0.16 ;
END MAS168

MACRO MAS169
   SIZE 0.08 BY 0.16 ;
END MAS169

MACRO MAS170
   SIZE 0.08 BY 0.16 ;
END MAS170

MACRO MAS171
   SIZE 0.08 BY 0.16 ;
END MAS171

MACRO MAS172
   SIZE 0.08 BY 0.16 ;
END MAS172

MACRO MAS173
   SIZE 0.08 BY 0.16 ;
END MAS173

MACRO MAS174
   SIZE 0.08 BY 0.16 ;
END MAS174

MACRO MAS175
   SIZE 0.08 BY 0.16 ;
END MAS175

MACRO MAS176
   SIZE 0.08 BY 0.16 ;
END MAS176

MACRO MAS177
   SIZE 0.08 BY 0.16 ;
END MAS177

MACRO MAS178
   SIZE 0.08 BY 0.16 ;
END MAS178

MACRO MAS179
   SIZE 0.08 BY 0.16 ;
END MAS179

MACRO MAS180
   SIZE 0.08 BY 0.16 ;
END MAS180

MACRO MAS181
   SIZE 0.08 BY 0.16 ;
END MAS181

MACRO MAS182
   SIZE 0.08 BY 0.16 ;
END MAS182

MACRO MAS183
   SIZE 0.08 BY 0.16 ;
END MAS183

MACRO MAS184
   SIZE 0.08 BY 0.16 ;
END MAS184

MACRO MAS185
   SIZE 0.08 BY 0.16 ;
END MAS185

MACRO MAS186
   SIZE 0.08 BY 0.16 ;
END MAS186

MACRO MAS187
   SIZE 0.08 BY 0.16 ;
END MAS187

MACRO MAS188
   SIZE 0.08 BY 0.16 ;
END MAS188

MACRO MAS189
   SIZE 0.08 BY 0.16 ;
END MAS189

MACRO MAS190
   SIZE 0.08 BY 0.16 ;
END MAS190

MACRO MAS191
   SIZE 0.08 BY 0.16 ;
END MAS191

MACRO MAS192
   SIZE 0.08 BY 0.16 ;
END MAS192

MACRO MAS193
   SIZE 0.08 BY 0.16 ;
END MAS193

MACRO MAS194
   SIZE 0.08 BY 0.16 ;
END MAS194

MACRO MAS195
   SIZE 0.08 BY 0.16 ;
END MAS195

MACRO MAS196
   SIZE 0.1 BY 0.16 ;
END MAS196

MACRO MAS197
   SIZE 0.1 BY 0.16 ;
END MAS197

MACRO MAS198
   SIZE 0.1 BY 0.16 ;
END MAS198

MACRO MAS199
   SIZE 0.1 BY 0.16 ;
END MAS199

MACRO MAS200
   SIZE 0.1 BY 0.16 ;
END MAS200

MACRO MAS201
   SIZE 0.1 BY 0.16 ;
END MAS201

MACRO MAS202
   SIZE 0.1 BY 0.16 ;
END MAS202

MACRO MAS203
   SIZE 0.1 BY 0.16 ;
END MAS203

MACRO MAS204
   SIZE 0.1 BY 0.16 ;
END MAS204

MACRO MAS205
   SIZE 0.1 BY 0.16 ;
END MAS205

MACRO MAS206
   SIZE 0.1 BY 0.16 ;
END MAS206

MACRO MAS207
   SIZE 0.1 BY 0.16 ;
END MAS207

MACRO MAS208
   SIZE 0.1 BY 0.16 ;
END MAS208

MACRO MAS209
   SIZE 0.1 BY 0.16 ;
END MAS209

MACRO MAS210
   SIZE 0.1 BY 0.16 ;
END MAS210

MACRO MAS211
   SIZE 0.1 BY 0.16 ;
END MAS211

MACRO MAS212
   SIZE 0.1 BY 0.16 ;
END MAS212

MACRO MAS213
   SIZE 0.1 BY 0.16 ;
END MAS213

MACRO MAS214
   SIZE 0.1 BY 0.16 ;
END MAS214

MACRO MAS215
   SIZE 0.1 BY 0.16 ;
END MAS215

MACRO MAS216
   SIZE 0.1 BY 0.16 ;
END MAS216

MACRO MAS217
   SIZE 0.1 BY 0.16 ;
END MAS217

MACRO MAS218
   SIZE 0.1 BY 0.16 ;
END MAS218

MACRO MAS219
   SIZE 0.1 BY 0.16 ;
END MAS219

MACRO MAS220
   SIZE 0.1 BY 0.16 ;
END MAS220

MACRO MAS221
   SIZE 0.1 BY 0.16 ;
END MAS221

MACRO MAS222
   SIZE 0.1 BY 0.16 ;
END MAS222

MACRO MAS223
   SIZE 0.1 BY 0.16 ;
END MAS223

MACRO MAS224
   SIZE 0.1 BY 0.16 ;
END MAS224

MACRO MAS225
   SIZE 0.1 BY 0.16 ;
END MAS225

MACRO MAS226
   SIZE 0.1 BY 0.16 ;
END MAS226

MACRO MAS227
   SIZE 0.1 BY 0.16 ;
END MAS227

MACRO MAS228
   SIZE 0.1 BY 0.16 ;
END MAS228

MACRO MAS229
   SIZE 0.1 BY 0.16 ;
END MAS229

MACRO MAS230
   SIZE 0.1 BY 0.16 ;
END MAS230

MACRO MAS231
   SIZE 0.1 BY 0.16 ;
END MAS231

MACRO MAS232
   SIZE 0.1 BY 0.16 ;
END MAS232

MACRO MAS233
   SIZE 0.1 BY 0.16 ;
END MAS233

MACRO MAS234
   SIZE 0.1 BY 0.16 ;
END MAS234

MACRO MAS235
   SIZE 0.1 BY 0.16 ;
END MAS235

MACRO MAS236
   SIZE 0.1 BY 0.16 ;
END MAS236

MACRO MAS237
   SIZE 0.1 BY 0.16 ;
END MAS237

MACRO MAS238
   SIZE 0.1 BY 0.16 ;
END MAS238

MACRO MAS239
   SIZE 0.1 BY 0.16 ;
END MAS239

MACRO MAS240
   SIZE 0.1 BY 0.16 ;
END MAS240

MACRO MAS241
   SIZE 0.1 BY 0.16 ;
END MAS241

MACRO MAS242
   SIZE 0.1 BY 0.16 ;
END MAS242

MACRO MAS243
   SIZE 0.1 BY 0.16 ;
END MAS243

MACRO MAS244
   SIZE 0.1 BY 0.16 ;
END MAS244

MACRO MAS245
   SIZE 0.1 BY 0.16 ;
END MAS245

MACRO MAS246
   SIZE 0.1 BY 0.16 ;
END MAS246

MACRO MAS247
   SIZE 0.1 BY 0.16 ;
END MAS247

MACRO MAS248
   SIZE 0.1 BY 0.16 ;
END MAS248

MACRO MAS249
   SIZE 0.1 BY 0.16 ;
END MAS249

MACRO MAS250
   SIZE 0.1 BY 0.16 ;
END MAS250

MACRO MAS251
   SIZE 0.1 BY 0.16 ;
END MAS251

MACRO MAS252
   SIZE 0.1 BY 0.16 ;
END MAS252

MACRO MAS253
   SIZE 0.1 BY 0.16 ;
END MAS253

MACRO MAS254
   SIZE 0.1 BY 0.16 ;
END MAS254

MACRO MAS255
   SIZE 0.1 BY 0.16 ;
END MAS255

MACRO MAS256
   SIZE 0.1 BY 0.16 ;
END MAS256

MACRO MAS257
   SIZE 0.1 BY 0.16 ;
END MAS257

MACRO MAS258
   SIZE 0.1 BY 0.16 ;
END MAS258

MACRO MAS259
   SIZE 0.1 BY 0.16 ;
END MAS259

MACRO MAS260
   SIZE 0.1 BY 0.16 ;
END MAS260

MACRO MAS261
   SIZE 0.1 BY 0.16 ;
END MAS261

MACRO MAS262
   SIZE 0.1 BY 0.16 ;
END MAS262

MACRO MAS263
   SIZE 0.1 BY 0.16 ;
END MAS263

MACRO MAS264
   SIZE 0.1 BY 0.16 ;
END MAS264

MACRO MAS265
   SIZE 0.1 BY 0.16 ;
END MAS265

MACRO MAS266
   SIZE 0.1 BY 0.16 ;
END MAS266

MACRO MAS267
   SIZE 0.1 BY 0.16 ;
END MAS267

MACRO MAS268
   SIZE 0.1 BY 0.16 ;
END MAS268

MACRO MAS269
   SIZE 0.1 BY 0.16 ;
END MAS269

MACRO MAS270
   SIZE 0.1 BY 0.16 ;
END MAS270

MACRO MAS271
   SIZE 0.1 BY 0.16 ;
END MAS271

MACRO MAS272
   SIZE 0.1 BY 0.16 ;
END MAS272

MACRO MAS273
   SIZE 0.1 BY 0.16 ;
END MAS273

MACRO MAS274
   SIZE 0.1 BY 0.16 ;
END MAS274

MACRO MAS275
   SIZE 0.1 BY 0.16 ;
END MAS275

MACRO MAS276
   SIZE 0.1 BY 0.16 ;
END MAS276

MACRO MAS277
   SIZE 0.1 BY 0.16 ;
END MAS277

MACRO MAS278
   SIZE 0.1 BY 0.16 ;
END MAS278

MACRO MAS279
   SIZE 0.1 BY 0.16 ;
END MAS279

MACRO MAS280
   SIZE 0.1 BY 0.16 ;
END MAS280

MACRO MAS281
   SIZE 0.1 BY 0.16 ;
END MAS281

MACRO MAS282
   SIZE 0.1 BY 0.16 ;
END MAS282

MACRO MAS283
   SIZE 0.1 BY 0.16 ;
END MAS283

MACRO MAS284
   SIZE 0.1 BY 0.16 ;
END MAS284

MACRO MAS285
   SIZE 0.1 BY 0.16 ;
END MAS285

MACRO MAS286
   SIZE 0.1 BY 0.16 ;
END MAS286

MACRO MAS287
   SIZE 0.1 BY 0.16 ;
END MAS287

MACRO MAS288
   SIZE 0.1 BY 0.16 ;
END MAS288

MACRO MAS289
   SIZE 0.1 BY 0.16 ;
END MAS289

MACRO MAS290
   SIZE 0.1 BY 0.16 ;
END MAS290

MACRO MAS291
   SIZE 0.1 BY 0.16 ;
END MAS291

MACRO MAS292
   SIZE 0.1 BY 0.16 ;
END MAS292

MACRO MAS293
   SIZE 0.1 BY 0.16 ;
END MAS293

MACRO MAS294
   SIZE 0.1 BY 0.16 ;
END MAS294

MACRO MAS295
   SIZE 0.1 BY 0.16 ;
END MAS295

MACRO MAS296
   SIZE 0.1 BY 0.16 ;
END MAS296

MACRO MAS297
   SIZE 0.1 BY 0.16 ;
END MAS297

MACRO MAS298
   SIZE 0.1 BY 0.16 ;
END MAS298

MACRO MAS299
   SIZE 0.1 BY 0.16 ;
END MAS299

MACRO MAS300
   SIZE 0.1 BY 0.16 ;
END MAS300

MACRO MAS301
   SIZE 0.1 BY 0.16 ;
END MAS301

MACRO MAS302
   SIZE 0.1 BY 0.16 ;
END MAS302

MACRO MAS303
   SIZE 0.1 BY 0.16 ;
END MAS303

MACRO MAS304
   SIZE 0.12 BY 0.16 ;
END MAS304

MACRO MAS305
   SIZE 0.12 BY 0.16 ;
END MAS305

MACRO MAS306
   SIZE 0.12 BY 0.16 ;
END MAS306

MACRO MAS307
   SIZE 0.12 BY 0.16 ;
END MAS307

MACRO MAS308
   SIZE 0.12 BY 0.16 ;
END MAS308

MACRO MAS309
   SIZE 0.12 BY 0.16 ;
END MAS309

MACRO MAS310
   SIZE 0.12 BY 0.16 ;
END MAS310

MACRO MAS311
   SIZE 0.12 BY 0.16 ;
END MAS311

MACRO MAS312
   SIZE 0.12 BY 0.16 ;
END MAS312

MACRO MAS313
   SIZE 0.12 BY 0.16 ;
END MAS313

MACRO MAS314
   SIZE 0.12 BY 0.16 ;
END MAS314

MACRO MAS315
   SIZE 0.12 BY 0.16 ;
END MAS315

MACRO MAS316
   SIZE 0.12 BY 0.16 ;
END MAS316

MACRO MAS317
   SIZE 0.12 BY 0.16 ;
END MAS317

MACRO MAS318
   SIZE 0.12 BY 0.16 ;
END MAS318

MACRO MAS319
   SIZE 0.12 BY 0.16 ;
END MAS319

MACRO MAS320
   SIZE 0.12 BY 0.16 ;
END MAS320

MACRO MAS321
   SIZE 0.12 BY 0.16 ;
END MAS321

MACRO MAS322
   SIZE 0.12 BY 0.16 ;
END MAS322

MACRO MAS323
   SIZE 0.12 BY 0.16 ;
END MAS323

MACRO MAS324
   SIZE 0.12 BY 0.16 ;
END MAS324

MACRO MAS325
   SIZE 0.12 BY 0.16 ;
END MAS325

MACRO MAS326
   SIZE 0.12 BY 0.16 ;
END MAS326

MACRO MAS327
   SIZE 0.12 BY 0.16 ;
END MAS327

MACRO MAS328
   SIZE 0.12 BY 0.16 ;
END MAS328

MACRO MAS329
   SIZE 0.12 BY 0.16 ;
END MAS329

MACRO MAS330
   SIZE 0.12 BY 0.16 ;
END MAS330

MACRO MAS331
   SIZE 0.12 BY 0.16 ;
END MAS331

MACRO MAS332
   SIZE 0.12 BY 0.16 ;
END MAS332

MACRO MAS333
   SIZE 0.12 BY 0.16 ;
END MAS333

MACRO MAS334
   SIZE 0.12 BY 0.16 ;
END MAS334

MACRO MAS335
   SIZE 0.12 BY 0.16 ;
END MAS335

MACRO MAS336
   SIZE 0.12 BY 0.16 ;
END MAS336

MACRO MAS337
   SIZE 0.12 BY 0.16 ;
END MAS337

MACRO MAS338
   SIZE 0.12 BY 0.16 ;
END MAS338

MACRO MAS339
   SIZE 0.12 BY 0.16 ;
END MAS339

MACRO MAS340
   SIZE 0.12 BY 0.16 ;
END MAS340

MACRO MAS341
   SIZE 0.12 BY 0.16 ;
END MAS341

MACRO MAS342
   SIZE 0.12 BY 0.16 ;
END MAS342

MACRO MAS343
   SIZE 0.12 BY 0.16 ;
END MAS343

MACRO MAS344
   SIZE 0.12 BY 0.16 ;
END MAS344

MACRO MAS345
   SIZE 0.12 BY 0.16 ;
END MAS345

MACRO MAS346
   SIZE 0.12 BY 0.16 ;
END MAS346

MACRO MAS347
   SIZE 0.12 BY 0.16 ;
END MAS347

MACRO MAS348
   SIZE 0.12 BY 0.16 ;
END MAS348

MACRO MAS349
   SIZE 0.12 BY 0.16 ;
END MAS349

MACRO MAS350
   SIZE 0.12 BY 0.16 ;
END MAS350

MACRO MAS351
   SIZE 0.12 BY 0.16 ;
END MAS351

MACRO MAS352
   SIZE 0.12 BY 0.16 ;
END MAS352

MACRO MAS353
   SIZE 0.12 BY 0.16 ;
END MAS353

MACRO MAS354
   SIZE 0.12 BY 0.16 ;
END MAS354

MACRO MAS355
   SIZE 0.12 BY 0.16 ;
END MAS355

MACRO MAS356
   SIZE 0.12 BY 0.16 ;
END MAS356

MACRO MAS357
   SIZE 0.12 BY 0.16 ;
END MAS357

MACRO MAS358
   SIZE 0.12 BY 0.16 ;
END MAS358

MACRO MAS359
   SIZE 0.12 BY 0.16 ;
END MAS359

MACRO MAS360
   SIZE 0.12 BY 0.16 ;
END MAS360

MACRO MAS361
   SIZE 0.12 BY 0.16 ;
END MAS361

MACRO MAS362
   SIZE 0.12 BY 0.16 ;
END MAS362

MACRO MAS363
   SIZE 0.12 BY 0.16 ;
END MAS363

MACRO MAS364
   SIZE 0.12 BY 0.16 ;
END MAS364

MACRO MAS365
   SIZE 0.12 BY 0.16 ;
END MAS365

MACRO MAS366
   SIZE 0.12 BY 0.16 ;
END MAS366

MACRO MAS367
   SIZE 0.12 BY 0.16 ;
END MAS367

MACRO MAS368
   SIZE 0.12 BY 0.16 ;
END MAS368

MACRO MAS369
   SIZE 0.12 BY 0.16 ;
END MAS369

MACRO MAS370
   SIZE 0.12 BY 0.16 ;
END MAS370

MACRO MAS371
   SIZE 0.12 BY 0.16 ;
END MAS371

MACRO MAS372
   SIZE 0.12 BY 0.16 ;
END MAS372

MACRO MAS373
   SIZE 0.12 BY 0.16 ;
END MAS373

MACRO MAS374
   SIZE 0.12 BY 0.16 ;
END MAS374

MACRO MAS375
   SIZE 0.12 BY 0.16 ;
END MAS375

MACRO MAS376
   SIZE 0.12 BY 0.16 ;
END MAS376

MACRO MAS377
   SIZE 0.12 BY 0.16 ;
END MAS377

MACRO MAS378
   SIZE 0.12 BY 0.16 ;
END MAS378

MACRO MAS379
   SIZE 0.12 BY 0.16 ;
END MAS379

MACRO MAS380
   SIZE 0.12 BY 0.16 ;
END MAS380

MACRO MAS381
   SIZE 0.12 BY 0.16 ;
END MAS381

MACRO MAS382
   SIZE 0.12 BY 0.16 ;
END MAS382

MACRO MAS383
   SIZE 0.12 BY 0.16 ;
END MAS383

MACRO MAS384
   SIZE 0.12 BY 0.16 ;
END MAS384

MACRO MAS385
   SIZE 0.12 BY 0.16 ;
END MAS385

MACRO MAS386
   SIZE 0.12 BY 0.16 ;
END MAS386

MACRO MAS387
   SIZE 0.12 BY 0.16 ;
END MAS387

MACRO MAS388
   SIZE 0.12 BY 0.16 ;
END MAS388

MACRO MAS389
   SIZE 0.12 BY 0.16 ;
END MAS389

MACRO MAS390
   SIZE 0.12 BY 0.16 ;
END MAS390

MACRO MAS391
   SIZE 0.12 BY 0.16 ;
END MAS391

MACRO MAS392
   SIZE 0.12 BY 0.16 ;
END MAS392

MACRO MAS393
   SIZE 0.12 BY 0.16 ;
END MAS393

MACRO MAS394
   SIZE 0.12 BY 0.16 ;
END MAS394

MACRO MAS395
   SIZE 0.12 BY 0.16 ;
END MAS395

MACRO MAS396
   SIZE 0.12 BY 0.16 ;
END MAS396

MACRO MAS397
   SIZE 0.12 BY 0.16 ;
END MAS397

MACRO MAS398
   SIZE 0.12 BY 0.16 ;
END MAS398

MACRO MAS399
   SIZE 0.12 BY 0.16 ;
END MAS399

MACRO MAS400
   SIZE 0.12 BY 0.16 ;
END MAS400

MACRO MAS401
   SIZE 0.12 BY 0.16 ;
END MAS401

MACRO MAS402
   SIZE 0.12 BY 0.16 ;
END MAS402

MACRO MAS403
   SIZE 0.12 BY 0.16 ;
END MAS403

MACRO MAS404
   SIZE 0.12 BY 0.16 ;
END MAS404

MACRO MAS405
   SIZE 0.12 BY 0.16 ;
END MAS405

MACRO MAS406
   SIZE 0.12 BY 0.16 ;
END MAS406

MACRO MAS407
   SIZE 0.12 BY 0.16 ;
END MAS407

MACRO MAS408
   SIZE 0.12 BY 0.16 ;
END MAS408

MACRO MAS409
   SIZE 0.12 BY 0.16 ;
END MAS409

MACRO MAS410
   SIZE 0.12 BY 0.16 ;
END MAS410

MACRO MAS411
   SIZE 0.12 BY 0.16 ;
END MAS411

MACRO MAS412
   SIZE 0.12 BY 0.16 ;
END MAS412

MACRO MAS413
   SIZE 0.12 BY 0.16 ;
END MAS413

MACRO MAS414
   SIZE 0.12 BY 0.16 ;
END MAS414

MACRO MAS415
   SIZE 0.12 BY 0.16 ;
END MAS415

MACRO MAS416
   SIZE 0.12 BY 0.16 ;
END MAS416

MACRO MAS417
   SIZE 0.12 BY 0.16 ;
END MAS417

MACRO MAS418
   SIZE 0.12 BY 0.16 ;
END MAS418

MACRO MAS419
   SIZE 0.12 BY 0.16 ;
END MAS419

MACRO MAS420
   SIZE 0.12 BY 0.16 ;
END MAS420

MACRO MAS421
   SIZE 0.12 BY 0.16 ;
END MAS421

MACRO MAS422
   SIZE 0.12 BY 0.16 ;
END MAS422

MACRO MAS423
   SIZE 0.12 BY 0.16 ;
END MAS423

MACRO MAS424
   SIZE 0.12 BY 0.16 ;
END MAS424

MACRO MAS425
   SIZE 0.12 BY 0.16 ;
END MAS425

MACRO MAS426
   SIZE 0.12 BY 0.16 ;
END MAS426

MACRO MAS427
   SIZE 0.12 BY 0.16 ;
END MAS427

MACRO MAS428
   SIZE 0.12 BY 0.16 ;
END MAS428

MACRO MAS429
   SIZE 0.12 BY 0.16 ;
END MAS429

MACRO MAS430
   SIZE 0.12 BY 0.16 ;
END MAS430

MACRO MAS431
   SIZE 0.12 BY 0.16 ;
END MAS431

MACRO MAS432
   SIZE 0.12 BY 0.16 ;
END MAS432

MACRO MAS433
   SIZE 0.12 BY 0.16 ;
END MAS433

MACRO MAS434
   SIZE 0.12 BY 0.16 ;
END MAS434

MACRO MAS435
   SIZE 0.12 BY 0.16 ;
END MAS435

MACRO MAS436
   SIZE 0.12 BY 0.16 ;
END MAS436

MACRO MAS437
   SIZE 0.12 BY 0.16 ;
END MAS437

MACRO MAS438
   SIZE 0.12 BY 0.16 ;
END MAS438

MACRO MAS439
   SIZE 0.12 BY 0.16 ;
END MAS439

MACRO MAS440
   SIZE 0.12 BY 0.16 ;
END MAS440

MACRO MAS441
   SIZE 0.12 BY 0.16 ;
END MAS441

MACRO MAS442
   SIZE 0.12 BY 0.16 ;
END MAS442

MACRO MAS443
   SIZE 0.12 BY 0.16 ;
END MAS443

MACRO MAS444
   SIZE 0.12 BY 0.16 ;
END MAS444

MACRO MAS445
   SIZE 0.12 BY 0.16 ;
END MAS445

MACRO MAS446
   SIZE 0.12 BY 0.16 ;
END MAS446

MACRO MAS447
   SIZE 0.12 BY 0.16 ;
END MAS447

MACRO MAS448
   SIZE 0.12 BY 0.16 ;
END MAS448

MACRO MAS449
   SIZE 0.12 BY 0.16 ;
END MAS449

MACRO MAS450
   SIZE 0.12 BY 0.16 ;
END MAS450

MACRO MAS451
   SIZE 0.12 BY 0.16 ;
END MAS451

MACRO MAS452
   SIZE 0.12 BY 0.16 ;
END MAS452

MACRO MAS453
   SIZE 0.12 BY 0.16 ;
END MAS453

MACRO MAS454
   SIZE 0.12 BY 0.16 ;
END MAS454

MACRO MAS455
   SIZE 0.12 BY 0.16 ;
END MAS455

MACRO MAS456
   SIZE 0.12 BY 0.16 ;
END MAS456

MACRO MAS457
   SIZE 0.12 BY 0.16 ;
END MAS457

MACRO MAS458
   SIZE 0.12 BY 0.16 ;
END MAS458

MACRO MAS459
   SIZE 0.12 BY 0.16 ;
END MAS459

MACRO MAS460
   SIZE 0.12 BY 0.16 ;
END MAS460

MACRO MAS461
   SIZE 0.12 BY 0.16 ;
END MAS461

MACRO MAS462
   SIZE 0.12 BY 0.16 ;
END MAS462

MACRO MAS463
   SIZE 0.12 BY 0.16 ;
END MAS463

MACRO MAS464
   SIZE 0.12 BY 0.16 ;
END MAS464

MACRO MAS465
   SIZE 0.12 BY 0.16 ;
END MAS465

MACRO MAS466
   SIZE 0.12 BY 0.16 ;
END MAS466

MACRO MAS467
   SIZE 0.12 BY 0.16 ;
END MAS467

MACRO MAS468
   SIZE 0.12 BY 0.16 ;
END MAS468

MACRO MAS469
   SIZE 0.12 BY 0.16 ;
END MAS469

MACRO MAS470
   SIZE 0.12 BY 0.16 ;
END MAS470

MACRO MAS471
   SIZE 0.12 BY 0.16 ;
END MAS471

MACRO MAS472
   SIZE 0.12 BY 0.16 ;
END MAS472

MACRO MAS473
   SIZE 0.12 BY 0.16 ;
END MAS473

MACRO MAS474
   SIZE 0.12 BY 0.16 ;
END MAS474

MACRO MAS475
   SIZE 0.12 BY 0.16 ;
END MAS475

MACRO MAS476
   SIZE 0.12 BY 0.16 ;
END MAS476

MACRO MAS477
   SIZE 0.12 BY 0.16 ;
END MAS477

MACRO MAS478
   SIZE 0.12 BY 0.16 ;
END MAS478

MACRO MAS479
   SIZE 0.12 BY 0.16 ;
END MAS479

MACRO MAS480
   SIZE 0.12 BY 0.16 ;
END MAS480

MACRO MAS481
   SIZE 0.12 BY 0.16 ;
END MAS481

MACRO MAS482
   SIZE 0.12 BY 0.16 ;
END MAS482

MACRO MAS483
   SIZE 0.12 BY 0.16 ;
END MAS483

MACRO MAS484
   SIZE 0.12 BY 0.16 ;
END MAS484

MACRO MAS485
   SIZE 0.12 BY 0.16 ;
END MAS485

MACRO MAS486
   SIZE 0.12 BY 0.16 ;
END MAS486

MACRO MAS487
   SIZE 0.12 BY 0.16 ;
END MAS487

MACRO MAS488
   SIZE 0.12 BY 0.16 ;
END MAS488

MACRO MAS489
   SIZE 0.12 BY 0.16 ;
END MAS489

MACRO MAS490
   SIZE 0.12 BY 0.16 ;
END MAS490

MACRO MAS491
   SIZE 0.12 BY 0.16 ;
END MAS491

MACRO MAS492
   SIZE 0.12 BY 0.16 ;
END MAS492

MACRO MAS493
   SIZE 0.12 BY 0.16 ;
END MAS493

MACRO MAS494
   SIZE 0.12 BY 0.16 ;
END MAS494

MACRO MAS495
   SIZE 0.12 BY 0.16 ;
END MAS495

MACRO MAS496
   SIZE 0.12 BY 0.16 ;
END MAS496

MACRO MAS497
   SIZE 0.12 BY 0.16 ;
END MAS497

MACRO MAS498
   SIZE 0.12 BY 0.16 ;
END MAS498

MACRO MAS499
   SIZE 0.12 BY 0.16 ;
END MAS499

MACRO MAS500
   SIZE 0.12 BY 0.16 ;
END MAS500

MACRO MAS501
   SIZE 0.12 BY 0.16 ;
END MAS501

MACRO MAS502
   SIZE 0.12 BY 0.16 ;
END MAS502

MACRO MAS503
   SIZE 0.12 BY 0.16 ;
END MAS503

MACRO MAS504
   SIZE 0.12 BY 0.16 ;
END MAS504

MACRO MAS505
   SIZE 0.12 BY 0.16 ;
END MAS505

MACRO MAS506
   SIZE 0.12 BY 0.16 ;
END MAS506

MACRO MAS507
   SIZE 0.12 BY 0.16 ;
END MAS507

MACRO MAS508
   SIZE 0.12 BY 0.16 ;
END MAS508

MACRO MAS509
   SIZE 0.12 BY 0.16 ;
END MAS509

MACRO MAS510
   SIZE 0.12 BY 0.16 ;
END MAS510

MACRO MAS511
   SIZE 0.12 BY 0.16 ;
END MAS511

MACRO MAS512
   SIZE 0.12 BY 0.16 ;
END MAS512

MACRO MAS513
   SIZE 0.12 BY 0.16 ;
END MAS513

MACRO MAS514
   SIZE 0.12 BY 0.16 ;
END MAS514

MACRO MAS515
   SIZE 0.12 BY 0.16 ;
END MAS515

MACRO MAS516
   SIZE 0.12 BY 0.16 ;
END MAS516

MACRO MAS517
   SIZE 0.12 BY 0.16 ;
END MAS517

MACRO MAS518
   SIZE 0.12 BY 0.16 ;
END MAS518

MACRO MAS519
   SIZE 0.12 BY 0.16 ;
END MAS519

MACRO MAS520
   SIZE 0.12 BY 0.16 ;
END MAS520

MACRO MAS521
   SIZE 0.12 BY 0.16 ;
END MAS521

MACRO MAS522
   SIZE 0.12 BY 0.16 ;
END MAS522

MACRO MAS523
   SIZE 0.12 BY 0.16 ;
END MAS523

MACRO MAS524
   SIZE 0.12 BY 0.16 ;
END MAS524

MACRO MAS525
   SIZE 0.12 BY 0.16 ;
END MAS525

MACRO MAS526
   SIZE 0.12 BY 0.16 ;
END MAS526

MACRO MAS527
   SIZE 0.12 BY 0.16 ;
END MAS527

MACRO MAS528
   SIZE 0.12 BY 0.16 ;
END MAS528

MACRO MAS529
   SIZE 0.12 BY 0.16 ;
END MAS529

MACRO MAS530
   SIZE 0.12 BY 0.16 ;
END MAS530

MACRO MAS531
   SIZE 0.12 BY 0.16 ;
END MAS531

MACRO MAS532
   SIZE 0.12 BY 0.16 ;
END MAS532

MACRO MAS533
   SIZE 0.12 BY 0.16 ;
END MAS533

MACRO MAS534
   SIZE 0.12 BY 0.16 ;
END MAS534

MACRO MAS535
   SIZE 0.12 BY 0.16 ;
END MAS535

MACRO MAS536
   SIZE 0.12 BY 0.16 ;
END MAS536

MACRO MAS537
   SIZE 0.12 BY 0.16 ;
END MAS537

MACRO MAS538
   SIZE 0.12 BY 0.16 ;
END MAS538

MACRO MAS539
   SIZE 0.12 BY 0.16 ;
END MAS539

MACRO MAS540
   SIZE 0.12 BY 0.16 ;
END MAS540

MACRO MAS541
   SIZE 0.12 BY 0.16 ;
END MAS541

MACRO MAS542
   SIZE 0.12 BY 0.16 ;
END MAS542

MACRO MAS543
   SIZE 0.12 BY 0.16 ;
END MAS543

MACRO MAS544
   SIZE 0.12 BY 0.16 ;
END MAS544

MACRO MAS545
   SIZE 0.12 BY 0.16 ;
END MAS545

MACRO MAS546
   SIZE 0.12 BY 0.16 ;
END MAS546

MACRO MAS547
   SIZE 0.12 BY 0.16 ;
END MAS547

MACRO MAS548
   SIZE 0.12 BY 0.16 ;
END MAS548

MACRO MAS549
   SIZE 0.12 BY 0.16 ;
END MAS549

MACRO MAS550
   SIZE 0.12 BY 0.16 ;
END MAS550

MACRO MAS551
   SIZE 0.12 BY 0.16 ;
END MAS551

MACRO MAS552
   SIZE 0.12 BY 0.16 ;
END MAS552

MACRO MAS553
   SIZE 0.12 BY 0.16 ;
END MAS553

MACRO MAS554
   SIZE 0.12 BY 0.16 ;
END MAS554

MACRO MAS555
   SIZE 0.12 BY 0.16 ;
END MAS555

MACRO MAS556
   SIZE 0.12 BY 0.16 ;
END MAS556

MACRO MAS557
   SIZE 0.12 BY 0.16 ;
END MAS557

MACRO MAS558
   SIZE 0.12 BY 0.16 ;
END MAS558

MACRO MAS559
   SIZE 0.12 BY 0.16 ;
END MAS559

MACRO MAS560
   SIZE 0.12 BY 0.16 ;
END MAS560

MACRO MAS561
   SIZE 0.12 BY 0.16 ;
END MAS561

MACRO MAS562
   SIZE 0.12 BY 0.16 ;
END MAS562

MACRO MAS563
   SIZE 0.12 BY 0.16 ;
END MAS563

MACRO MAS564
   SIZE 0.12 BY 0.16 ;
END MAS564

MACRO MAS565
   SIZE 0.12 BY 0.16 ;
END MAS565

MACRO MAS566
   SIZE 0.12 BY 0.16 ;
END MAS566

MACRO MAS567
   SIZE 0.12 BY 0.16 ;
END MAS567

MACRO MAS568
   SIZE 0.12 BY 0.16 ;
END MAS568

MACRO MAS569
   SIZE 0.12 BY 0.16 ;
END MAS569

MACRO MAS570
   SIZE 0.12 BY 0.16 ;
END MAS570

MACRO MAS571
   SIZE 0.12 BY 0.16 ;
END MAS571

MACRO MAS572
   SIZE 0.12 BY 0.16 ;
END MAS572

MACRO MAS573
   SIZE 0.12 BY 0.16 ;
END MAS573

MACRO MAS574
   SIZE 0.12 BY 0.16 ;
END MAS574

MACRO MAS575
   SIZE 0.12 BY 0.16 ;
END MAS575

MACRO MAS576
   SIZE 0.12 BY 0.16 ;
END MAS576

MACRO MAS577
   SIZE 0.12 BY 0.16 ;
END MAS577

MACRO MAS578
   SIZE 0.12 BY 0.16 ;
END MAS578

MACRO MAS579
   SIZE 0.12 BY 0.16 ;
END MAS579

MACRO MAS580
   SIZE 0.12 BY 0.16 ;
END MAS580

MACRO MAS581
   SIZE 0.12 BY 0.16 ;
END MAS581

MACRO MAS582
   SIZE 0.12 BY 0.16 ;
END MAS582

MACRO MAS583
   SIZE 0.12 BY 0.16 ;
END MAS583

MACRO MAS584
   SIZE 0.12 BY 0.16 ;
END MAS584

MACRO MAS585
   SIZE 0.12 BY 0.16 ;
END MAS585

MACRO MAS586
   SIZE 0.12 BY 0.16 ;
END MAS586

MACRO MAS587
   SIZE 0.12 BY 0.16 ;
END MAS587

MACRO MAS588
   SIZE 0.12 BY 0.16 ;
END MAS588

MACRO MAS589
   SIZE 0.12 BY 0.16 ;
END MAS589

MACRO MAS590
   SIZE 0.12 BY 0.16 ;
END MAS590

MACRO MAS591
   SIZE 0.12 BY 0.16 ;
END MAS591

MACRO MAS592
   SIZE 0.12 BY 0.16 ;
END MAS592

MACRO MAS593
   SIZE 0.12 BY 0.16 ;
END MAS593

MACRO MAS594
   SIZE 0.12 BY 0.16 ;
END MAS594

MACRO MAS595
   SIZE 0.12 BY 0.16 ;
END MAS595

MACRO MAS596
   SIZE 0.12 BY 0.16 ;
END MAS596

MACRO MAS597
   SIZE 0.12 BY 0.16 ;
END MAS597

MACRO MAS598
   SIZE 0.12 BY 0.16 ;
END MAS598

MACRO MAS599
   SIZE 0.12 BY 0.16 ;
END MAS599

MACRO MAS600
   SIZE 0.12 BY 0.16 ;
END MAS600

MACRO MAS601
   SIZE 0.12 BY 0.16 ;
END MAS601

MACRO MAS602
   SIZE 0.12 BY 0.16 ;
END MAS602

MACRO MAS603
   SIZE 0.12 BY 0.16 ;
END MAS603

MACRO MAS604
   SIZE 0.12 BY 0.16 ;
END MAS604

MACRO MAS605
   SIZE 0.12 BY 0.16 ;
END MAS605

MACRO MAS606
   SIZE 0.12 BY 0.16 ;
END MAS606

MACRO MAS607
   SIZE 0.12 BY 0.16 ;
END MAS607

MACRO MAS608
   SIZE 0.12 BY 0.16 ;
END MAS608

MACRO MAS609
   SIZE 0.12 BY 0.16 ;
END MAS609

MACRO MAS610
   SIZE 0.12 BY 0.16 ;
END MAS610

MACRO MAS611
   SIZE 0.12 BY 0.16 ;
END MAS611

MACRO MAS612
   SIZE 0.12 BY 0.16 ;
END MAS612

MACRO MAS613
   SIZE 0.12 BY 0.16 ;
END MAS613

MACRO MAS614
   SIZE 0.12 BY 0.16 ;
END MAS614

MACRO MAS615
   SIZE 0.12 BY 0.16 ;
END MAS615

MACRO MAS616
   SIZE 0.12 BY 0.16 ;
END MAS616

MACRO MAS617
   SIZE 0.12 BY 0.16 ;
END MAS617

MACRO MAS618
   SIZE 0.12 BY 0.16 ;
END MAS618

MACRO MAS619
   SIZE 0.12 BY 0.16 ;
END MAS619

MACRO MAS620
   SIZE 0.12 BY 0.16 ;
END MAS620

MACRO MAS621
   SIZE 0.12 BY 0.16 ;
END MAS621

MACRO MAS622
   SIZE 0.12 BY 0.16 ;
END MAS622

MACRO MAS623
   SIZE 0.12 BY 0.16 ;
END MAS623

MACRO MAS624
   SIZE 0.12 BY 0.16 ;
END MAS624

MACRO MAS625
   SIZE 0.12 BY 0.16 ;
END MAS625

MACRO MAS626
   SIZE 0.12 BY 0.16 ;
END MAS626

MACRO MAS627
   SIZE 0.12 BY 0.16 ;
END MAS627

MACRO MAS628
   SIZE 0.12 BY 0.16 ;
END MAS628

MACRO MAS629
   SIZE 0.12 BY 0.16 ;
END MAS629

MACRO MAS630
   SIZE 0.12 BY 0.16 ;
END MAS630

MACRO MAS631
   SIZE 0.12 BY 0.16 ;
END MAS631

MACRO MAS632
   SIZE 0.12 BY 0.16 ;
END MAS632

MACRO MAS633
   SIZE 0.12 BY 0.16 ;
END MAS633

MACRO MAS634
   SIZE 0.12 BY 0.16 ;
END MAS634

MACRO MAS635
   SIZE 0.12 BY 0.16 ;
END MAS635

MACRO MAS636
   SIZE 0.12 BY 0.16 ;
END MAS636

MACRO MAS637
   SIZE 0.12 BY 0.16 ;
END MAS637

MACRO MAS638
   SIZE 0.12 BY 0.16 ;
END MAS638

MACRO MAS639
   SIZE 0.12 BY 0.16 ;
END MAS639

MACRO MAS640
   SIZE 0.12 BY 0.16 ;
END MAS640

MACRO MAS641
   SIZE 0.12 BY 0.16 ;
END MAS641

MACRO MAS642
   SIZE 0.12 BY 0.16 ;
END MAS642

MACRO MAS643
   SIZE 0.12 BY 0.16 ;
END MAS643

MACRO MAS644
   SIZE 0.12 BY 0.16 ;
END MAS644

MACRO MAS645
   SIZE 0.12 BY 0.16 ;
END MAS645

MACRO MAS646
   SIZE 0.12 BY 0.16 ;
END MAS646

MACRO MAS647
   SIZE 0.12 BY 0.16 ;
END MAS647

MACRO MAS648
   SIZE 0.12 BY 0.16 ;
END MAS648

MACRO MAS649
   SIZE 0.12 BY 0.16 ;
END MAS649

MACRO MAS650
   SIZE 0.12 BY 0.16 ;
END MAS650

MACRO MAS651
   SIZE 0.12 BY 0.16 ;
END MAS651

MACRO MAS652
   SIZE 0.12 BY 0.16 ;
END MAS652

MACRO MAS653
   SIZE 0.12 BY 0.16 ;
END MAS653

MACRO MAS654
   SIZE 0.12 BY 0.16 ;
END MAS654

MACRO MAS655
   SIZE 0.12 BY 0.16 ;
END MAS655

MACRO MAS656
   SIZE 0.12 BY 0.16 ;
END MAS656

MACRO MAS657
   SIZE 0.12 BY 0.16 ;
END MAS657

MACRO MAS658
   SIZE 0.12 BY 0.16 ;
END MAS658

MACRO MAS659
   SIZE 0.12 BY 0.16 ;
END MAS659

MACRO MAS660
   SIZE 0.12 BY 0.16 ;
END MAS660

MACRO MAS661
   SIZE 0.12 BY 0.16 ;
END MAS661

MACRO MAS662
   SIZE 0.12 BY 0.16 ;
END MAS662

MACRO MAS663
   SIZE 0.12 BY 0.16 ;
END MAS663

MACRO MAS664
   SIZE 0.12 BY 0.16 ;
END MAS664

MACRO MAS665
   SIZE 0.12 BY 0.16 ;
END MAS665

MACRO MAS666
   SIZE 0.12 BY 0.16 ;
END MAS666

MACRO MAS667
   SIZE 0.12 BY 0.16 ;
END MAS667

MACRO MAS668
   SIZE 0.12 BY 0.16 ;
END MAS668

MACRO MAS669
   SIZE 0.12 BY 0.16 ;
END MAS669

MACRO MAS670
   SIZE 0.12 BY 0.16 ;
END MAS670

MACRO MAS671
   SIZE 0.12 BY 0.16 ;
END MAS671

MACRO MAS672
   SIZE 0.12 BY 0.16 ;
END MAS672

MACRO MAS673
   SIZE 0.12 BY 0.16 ;
END MAS673

MACRO MAS674
   SIZE 0.12 BY 0.16 ;
END MAS674

MACRO MAS675
   SIZE 0.12 BY 0.16 ;
END MAS675

MACRO MAS676
   SIZE 0.12 BY 0.16 ;
END MAS676

MACRO MAS677
   SIZE 0.12 BY 0.16 ;
END MAS677

MACRO MAS678
   SIZE 0.12 BY 0.16 ;
END MAS678

MACRO MAS679
   SIZE 0.12 BY 0.16 ;
END MAS679

MACRO MAS680
   SIZE 0.12 BY 0.16 ;
END MAS680

MACRO MAS681
   SIZE 0.12 BY 0.16 ;
END MAS681

MACRO MAS682
   SIZE 0.12 BY 0.16 ;
END MAS682

MACRO MAS683
   SIZE 0.12 BY 0.16 ;
END MAS683

MACRO MAS684
   SIZE 0.12 BY 0.16 ;
END MAS684

MACRO MAS685
   SIZE 0.12 BY 0.16 ;
END MAS685

MACRO MAS686
   SIZE 0.12 BY 0.16 ;
END MAS686

MACRO MAS687
   SIZE 0.12 BY 0.16 ;
END MAS687

MACRO MAS688
   SIZE 0.12 BY 0.16 ;
END MAS688

MACRO MAS689
   SIZE 0.12 BY 0.16 ;
END MAS689

MACRO MAS690
   SIZE 0.12 BY 0.16 ;
END MAS690

MACRO MAS691
   SIZE 0.12 BY 0.16 ;
END MAS691

MACRO MAS692
   SIZE 0.12 BY 0.16 ;
END MAS692

MACRO MAS693
   SIZE 0.12 BY 0.16 ;
END MAS693

MACRO MAS694
   SIZE 0.12 BY 0.16 ;
END MAS694

MACRO MAS695
   SIZE 0.12 BY 0.16 ;
END MAS695

MACRO MAS696
   SIZE 0.12 BY 0.16 ;
END MAS696

MACRO MAS697
   SIZE 0.12 BY 0.16 ;
END MAS697

MACRO MAS698
   SIZE 0.14 BY 0.16 ;
END MAS698

MACRO MAS699
   SIZE 0.14 BY 0.16 ;
END MAS699

MACRO MAS700
   SIZE 0.14 BY 0.16 ;
END MAS700

MACRO MAS701
   SIZE 0.14 BY 0.16 ;
END MAS701

MACRO MAS702
   SIZE 0.14 BY 0.16 ;
END MAS702

MACRO MAS703
   SIZE 0.14 BY 0.16 ;
END MAS703

MACRO MAS704
   SIZE 0.14 BY 0.16 ;
END MAS704

MACRO MAS705
   SIZE 0.14 BY 0.16 ;
END MAS705

MACRO MAS706
   SIZE 0.14 BY 0.16 ;
END MAS706

MACRO MAS707
   SIZE 0.14 BY 0.16 ;
END MAS707

MACRO MAS708
   SIZE 0.14 BY 0.16 ;
END MAS708

MACRO MAS709
   SIZE 0.14 BY 0.16 ;
END MAS709

MACRO MAS710
   SIZE 0.14 BY 0.16 ;
END MAS710

MACRO MAS711
   SIZE 0.14 BY 0.16 ;
END MAS711

MACRO MAS712
   SIZE 0.14 BY 0.16 ;
END MAS712

MACRO MAS713
   SIZE 0.14 BY 0.16 ;
END MAS713

MACRO MAS714
   SIZE 0.14 BY 0.16 ;
END MAS714

MACRO MAS715
   SIZE 0.14 BY 0.16 ;
END MAS715

MACRO MAS716
   SIZE 0.14 BY 0.16 ;
END MAS716

MACRO MAS717
   SIZE 0.14 BY 0.16 ;
END MAS717

MACRO MAS718
   SIZE 0.14 BY 0.16 ;
END MAS718

MACRO MAS719
   SIZE 0.14 BY 0.16 ;
END MAS719

MACRO MAS720
   SIZE 0.14 BY 0.16 ;
END MAS720

MACRO MAS721
   SIZE 0.14 BY 0.16 ;
END MAS721

MACRO MAS722
   SIZE 0.14 BY 0.16 ;
END MAS722

MACRO MAS723
   SIZE 0.14 BY 0.16 ;
END MAS723

MACRO MAS724
   SIZE 0.14 BY 0.16 ;
END MAS724

MACRO MAS725
   SIZE 0.14 BY 0.16 ;
END MAS725

MACRO MAS726
   SIZE 0.14 BY 0.16 ;
END MAS726

MACRO MAS727
   SIZE 0.14 BY 0.16 ;
END MAS727

MACRO MAS728
   SIZE 0.14 BY 0.16 ;
END MAS728

MACRO MAS729
   SIZE 0.14 BY 0.16 ;
END MAS729

MACRO MAS730
   SIZE 0.14 BY 0.16 ;
END MAS730

MACRO MAS731
   SIZE 0.14 BY 0.16 ;
END MAS731

MACRO MAS732
   SIZE 0.14 BY 0.16 ;
END MAS732

MACRO MAS733
   SIZE 0.14 BY 0.16 ;
END MAS733

MACRO MAS734
   SIZE 0.14 BY 0.16 ;
END MAS734

MACRO MAS735
   SIZE 0.14 BY 0.16 ;
END MAS735

MACRO MAS736
   SIZE 0.14 BY 0.16 ;
END MAS736

MACRO MAS737
   SIZE 0.14 BY 0.16 ;
END MAS737

MACRO MAS738
   SIZE 0.14 BY 0.16 ;
END MAS738

MACRO MAS739
   SIZE 0.14 BY 0.16 ;
END MAS739

MACRO MAS740
   SIZE 0.14 BY 0.16 ;
END MAS740

MACRO MAS741
   SIZE 0.14 BY 0.16 ;
END MAS741

MACRO MAS742
   SIZE 0.14 BY 0.16 ;
END MAS742

MACRO MAS743
   SIZE 0.14 BY 0.16 ;
END MAS743

MACRO MAS744
   SIZE 0.14 BY 0.16 ;
END MAS744

MACRO MAS745
   SIZE 0.14 BY 0.16 ;
END MAS745

MACRO MAS746
   SIZE 0.14 BY 0.16 ;
END MAS746

MACRO MAS747
   SIZE 0.14 BY 0.16 ;
END MAS747

MACRO MAS748
   SIZE 0.14 BY 0.16 ;
END MAS748

MACRO MAS749
   SIZE 0.14 BY 0.16 ;
END MAS749

MACRO MAS750
   SIZE 0.14 BY 0.16 ;
END MAS750

MACRO MAS751
   SIZE 0.14 BY 0.16 ;
END MAS751

MACRO MAS752
   SIZE 0.14 BY 0.16 ;
END MAS752

MACRO MAS753
   SIZE 0.14 BY 0.16 ;
END MAS753

MACRO MAS754
   SIZE 0.14 BY 0.16 ;
END MAS754

MACRO MAS755
   SIZE 0.14 BY 0.16 ;
END MAS755

MACRO MAS756
   SIZE 0.14 BY 0.16 ;
END MAS756

MACRO MAS757
   SIZE 0.14 BY 0.16 ;
END MAS757

MACRO MAS758
   SIZE 0.14 BY 0.16 ;
END MAS758

MACRO MAS759
   SIZE 0.14 BY 0.16 ;
END MAS759

MACRO MAS760
   SIZE 0.14 BY 0.16 ;
END MAS760

MACRO MAS761
   SIZE 0.14 BY 0.16 ;
END MAS761

MACRO MAS762
   SIZE 0.14 BY 0.16 ;
END MAS762

MACRO MAS763
   SIZE 0.14 BY 0.16 ;
END MAS763

MACRO MAS764
   SIZE 0.14 BY 0.16 ;
END MAS764

MACRO MAS765
   SIZE 0.14 BY 0.16 ;
END MAS765

MACRO MAS766
   SIZE 0.14 BY 0.16 ;
END MAS766

MACRO MAS767
   SIZE 0.14 BY 0.16 ;
END MAS767

MACRO MAS768
   SIZE 0.14 BY 0.16 ;
END MAS768

MACRO MAS769
   SIZE 0.14 BY 0.16 ;
END MAS769

MACRO MAS770
   SIZE 0.14 BY 0.16 ;
END MAS770

MACRO MAS771
   SIZE 0.14 BY 0.16 ;
END MAS771

MACRO MAS772
   SIZE 0.14 BY 0.16 ;
END MAS772

MACRO MAS773
   SIZE 0.14 BY 0.16 ;
END MAS773

MACRO MAS774
   SIZE 0.14 BY 0.16 ;
END MAS774

MACRO MAS775
   SIZE 0.14 BY 0.16 ;
END MAS775

MACRO MAS776
   SIZE 0.14 BY 0.16 ;
END MAS776

MACRO MAS777
   SIZE 0.14 BY 0.16 ;
END MAS777

MACRO MAS778
   SIZE 0.14 BY 0.16 ;
END MAS778

MACRO MAS779
   SIZE 0.14 BY 0.16 ;
END MAS779

MACRO MAS780
   SIZE 0.14 BY 0.16 ;
END MAS780

MACRO MAS781
   SIZE 0.14 BY 0.16 ;
END MAS781

MACRO MAS782
   SIZE 0.14 BY 0.16 ;
END MAS782

MACRO MAS783
   SIZE 0.14 BY 0.16 ;
END MAS783

MACRO MAS784
   SIZE 0.14 BY 0.16 ;
END MAS784

MACRO MAS785
   SIZE 0.14 BY 0.16 ;
END MAS785

MACRO MAS786
   SIZE 0.14 BY 0.16 ;
END MAS786

MACRO MAS787
   SIZE 0.14 BY 0.16 ;
END MAS787

MACRO MAS788
   SIZE 0.14 BY 0.16 ;
END MAS788

MACRO MAS789
   SIZE 0.14 BY 0.16 ;
END MAS789

MACRO MAS790
   SIZE 0.14 BY 0.16 ;
END MAS790

MACRO MAS791
   SIZE 0.14 BY 0.16 ;
END MAS791

MACRO MAS792
   SIZE 0.14 BY 0.16 ;
END MAS792

MACRO MAS793
   SIZE 0.14 BY 0.16 ;
END MAS793

MACRO MAS794
   SIZE 0.14 BY 0.16 ;
END MAS794

MACRO MAS795
   SIZE 0.14 BY 0.16 ;
END MAS795

MACRO MAS796
   SIZE 0.14 BY 0.16 ;
END MAS796

MACRO MAS797
   SIZE 0.14 BY 0.16 ;
END MAS797

MACRO MAS798
   SIZE 0.14 BY 0.16 ;
END MAS798

MACRO MAS799
   SIZE 0.14 BY 0.16 ;
END MAS799

MACRO MAS800
   SIZE 0.14 BY 0.16 ;
END MAS800

MACRO MAS801
   SIZE 0.14 BY 0.16 ;
END MAS801

MACRO MAS802
   SIZE 0.14 BY 0.16 ;
END MAS802

MACRO MAS803
   SIZE 0.14 BY 0.16 ;
END MAS803

MACRO MAS804
   SIZE 0.14 BY 0.16 ;
END MAS804

MACRO MAS805
   SIZE 0.14 BY 0.16 ;
END MAS805

MACRO MAS806
   SIZE 0.14 BY 0.16 ;
END MAS806

MACRO MAS807
   SIZE 0.14 BY 0.16 ;
END MAS807

MACRO MAS808
   SIZE 0.14 BY 0.16 ;
END MAS808

MACRO MAS809
   SIZE 0.14 BY 0.16 ;
END MAS809

MACRO MAS810
   SIZE 0.14 BY 0.16 ;
END MAS810

MACRO MAS811
   SIZE 0.14 BY 0.16 ;
END MAS811

MACRO MAS812
   SIZE 0.14 BY 0.16 ;
END MAS812

MACRO MAS813
   SIZE 0.14 BY 0.16 ;
END MAS813

MACRO MAS814
   SIZE 0.14 BY 0.16 ;
END MAS814

MACRO MAS815
   SIZE 0.14 BY 0.16 ;
END MAS815

MACRO MAS816
   SIZE 0.14 BY 0.16 ;
END MAS816

MACRO MAS817
   SIZE 0.14 BY 0.16 ;
END MAS817

MACRO MAS818
   SIZE 0.14 BY 0.16 ;
END MAS818

MACRO MAS819
   SIZE 0.14 BY 0.16 ;
END MAS819

MACRO MAS820
   SIZE 0.14 BY 0.16 ;
END MAS820

MACRO MAS821
   SIZE 0.14 BY 0.16 ;
END MAS821

MACRO MAS822
   SIZE 0.14 BY 0.16 ;
END MAS822

MACRO MAS823
   SIZE 0.14 BY 0.16 ;
END MAS823

MACRO MAS824
   SIZE 0.14 BY 0.16 ;
END MAS824

MACRO MAS825
   SIZE 0.14 BY 0.16 ;
END MAS825

MACRO MAS826
   SIZE 0.14 BY 0.16 ;
END MAS826

MACRO MAS827
   SIZE 0.14 BY 0.16 ;
END MAS827

MACRO MAS828
   SIZE 0.14 BY 0.16 ;
END MAS828

MACRO MAS829
   SIZE 0.14 BY 0.16 ;
END MAS829

MACRO MAS830
   SIZE 0.14 BY 0.16 ;
END MAS830

MACRO MAS831
   SIZE 0.14 BY 0.16 ;
END MAS831

MACRO MAS832
   SIZE 0.14 BY 0.16 ;
END MAS832

MACRO MAS833
   SIZE 0.14 BY 0.16 ;
END MAS833

MACRO MAS834
   SIZE 0.14 BY 0.16 ;
END MAS834

MACRO MAS835
   SIZE 0.14 BY 0.16 ;
END MAS835

MACRO MAS836
   SIZE 0.14 BY 0.16 ;
END MAS836

MACRO MAS837
   SIZE 0.14 BY 0.16 ;
END MAS837

MACRO MAS838
   SIZE 0.14 BY 0.16 ;
END MAS838

MACRO MAS839
   SIZE 0.14 BY 0.16 ;
END MAS839

MACRO MAS840
   SIZE 0.14 BY 0.16 ;
END MAS840

MACRO MAS841
   SIZE 0.14 BY 0.16 ;
END MAS841

MACRO MAS842
   SIZE 0.14 BY 0.16 ;
END MAS842

MACRO MAS843
   SIZE 0.14 BY 0.16 ;
END MAS843

MACRO MAS844
   SIZE 0.14 BY 0.16 ;
END MAS844

MACRO MAS845
   SIZE 0.14 BY 0.16 ;
END MAS845

MACRO MAS846
   SIZE 0.14 BY 0.16 ;
END MAS846

MACRO MAS847
   SIZE 0.14 BY 0.16 ;
END MAS847

MACRO MAS848
   SIZE 0.14 BY 0.16 ;
END MAS848

MACRO MAS849
   SIZE 0.14 BY 0.16 ;
END MAS849

MACRO MAS850
   SIZE 0.14 BY 0.16 ;
END MAS850

MACRO MAS851
   SIZE 0.14 BY 0.16 ;
END MAS851

MACRO MAS852
   SIZE 0.14 BY 0.16 ;
END MAS852

MACRO MAS853
   SIZE 0.14 BY 0.16 ;
END MAS853

MACRO MAS854
   SIZE 0.14 BY 0.16 ;
END MAS854

MACRO MAS855
   SIZE 0.14 BY 0.16 ;
END MAS855

MACRO MAS856
   SIZE 0.14 BY 0.16 ;
END MAS856

MACRO MAS857
   SIZE 0.14 BY 0.16 ;
END MAS857

MACRO MAS858
   SIZE 0.14 BY 0.16 ;
END MAS858

MACRO MAS859
   SIZE 0.14 BY 0.16 ;
END MAS859

MACRO MAS860
   SIZE 0.14 BY 0.16 ;
END MAS860

MACRO MAS861
   SIZE 0.14 BY 0.16 ;
END MAS861

MACRO MAS862
   SIZE 0.14 BY 0.16 ;
END MAS862

MACRO MAS863
   SIZE 0.14 BY 0.16 ;
END MAS863

MACRO MAS864
   SIZE 0.14 BY 0.16 ;
END MAS864

MACRO MAS865
   SIZE 0.14 BY 0.16 ;
END MAS865

MACRO MAS866
   SIZE 0.14 BY 0.16 ;
END MAS866

MACRO MAS867
   SIZE 0.14 BY 0.16 ;
END MAS867

MACRO MAS868
   SIZE 0.14 BY 0.16 ;
END MAS868

MACRO MAS869
   SIZE 0.14 BY 0.16 ;
END MAS869

MACRO MAS870
   SIZE 0.14 BY 0.16 ;
END MAS870

MACRO MAS871
   SIZE 0.14 BY 0.16 ;
END MAS871

MACRO MAS872
   SIZE 0.14 BY 0.16 ;
END MAS872

MACRO MAS873
   SIZE 0.14 BY 0.16 ;
END MAS873

MACRO MAS874
   SIZE 0.14 BY 0.16 ;
END MAS874

MACRO MAS875
   SIZE 0.14 BY 0.16 ;
END MAS875

MACRO MAS876
   SIZE 0.14 BY 0.16 ;
END MAS876

MACRO MAS877
   SIZE 0.14 BY 0.16 ;
END MAS877

MACRO MAS878
   SIZE 0.14 BY 0.16 ;
END MAS878

MACRO MAS879
   SIZE 0.14 BY 0.16 ;
END MAS879

MACRO MAS880
   SIZE 0.14 BY 0.16 ;
END MAS880

MACRO MAS881
   SIZE 0.14 BY 0.16 ;
END MAS881

MACRO MAS882
   SIZE 0.14 BY 0.16 ;
END MAS882

MACRO MAS883
   SIZE 0.14 BY 0.16 ;
END MAS883

MACRO MAS884
   SIZE 0.14 BY 0.16 ;
END MAS884

MACRO MAS885
   SIZE 0.14 BY 0.16 ;
END MAS885

MACRO MAS886
   SIZE 0.14 BY 0.16 ;
END MAS886

MACRO MAS887
   SIZE 0.14 BY 0.16 ;
END MAS887

MACRO MAS888
   SIZE 0.14 BY 0.16 ;
END MAS888

MACRO MAS889
   SIZE 0.14 BY 0.16 ;
END MAS889

MACRO MAS890
   SIZE 0.14 BY 0.16 ;
END MAS890

MACRO MAS891
   SIZE 0.14 BY 0.16 ;
END MAS891

MACRO MAS892
   SIZE 0.14 BY 0.16 ;
END MAS892

MACRO MAS893
   SIZE 0.14 BY 0.16 ;
END MAS893

MACRO MAS894
   SIZE 0.14 BY 0.16 ;
END MAS894

MACRO MAS895
   SIZE 0.14 BY 0.16 ;
END MAS895

MACRO MAS896
   SIZE 0.14 BY 0.16 ;
END MAS896

MACRO MAS897
   SIZE 0.14 BY 0.16 ;
END MAS897

MACRO MAS898
   SIZE 0.14 BY 0.16 ;
END MAS898

MACRO MAS899
   SIZE 0.14 BY 0.16 ;
END MAS899

MACRO MAS900
   SIZE 0.14 BY 0.16 ;
END MAS900

MACRO MAS901
   SIZE 0.14 BY 0.16 ;
END MAS901

MACRO MAS902
   SIZE 0.14 BY 0.16 ;
END MAS902

MACRO MAS903
   SIZE 0.14 BY 0.16 ;
END MAS903

MACRO MAS904
   SIZE 0.14 BY 0.16 ;
END MAS904

MACRO MAS905
   SIZE 0.14 BY 0.16 ;
END MAS905

MACRO MAS906
   SIZE 0.14 BY 0.16 ;
END MAS906

MACRO MAS907
   SIZE 0.14 BY 0.16 ;
END MAS907

MACRO MAS908
   SIZE 0.14 BY 0.16 ;
END MAS908

MACRO MAS909
   SIZE 0.14 BY 0.16 ;
END MAS909

MACRO MAS910
   SIZE 0.14 BY 0.16 ;
END MAS910

MACRO MAS911
   SIZE 0.14 BY 0.16 ;
END MAS911

MACRO MAS912
   SIZE 0.14 BY 0.16 ;
END MAS912

MACRO MAS913
   SIZE 0.14 BY 0.16 ;
END MAS913

MACRO MAS914
   SIZE 0.14 BY 0.16 ;
END MAS914

MACRO MAS915
   SIZE 0.14 BY 0.16 ;
END MAS915

MACRO MAS916
   SIZE 0.14 BY 0.16 ;
END MAS916

MACRO MAS917
   SIZE 0.14 BY 0.16 ;
END MAS917

MACRO MAS918
   SIZE 0.14 BY 0.16 ;
END MAS918

MACRO MAS919
   SIZE 0.14 BY 0.16 ;
END MAS919

MACRO MAS920
   SIZE 0.14 BY 0.16 ;
END MAS920

MACRO MAS921
   SIZE 0.14 BY 0.16 ;
END MAS921

MACRO MAS922
   SIZE 0.14 BY 0.16 ;
END MAS922

MACRO MAS923
   SIZE 0.14 BY 0.16 ;
END MAS923

MACRO MAS924
   SIZE 0.14 BY 0.16 ;
END MAS924

MACRO MAS925
   SIZE 0.14 BY 0.16 ;
END MAS925

MACRO MAS926
   SIZE 0.14 BY 0.16 ;
END MAS926

MACRO MAS927
   SIZE 0.14 BY 0.16 ;
END MAS927

MACRO MAS928
   SIZE 0.14 BY 0.16 ;
END MAS928

MACRO MAS929
   SIZE 0.14 BY 0.16 ;
END MAS929

MACRO MAS930
   SIZE 0.14 BY 0.16 ;
END MAS930

MACRO MAS931
   SIZE 0.14 BY 0.16 ;
END MAS931

MACRO MAS932
   SIZE 0.14 BY 0.16 ;
END MAS932

MACRO MAS933
   SIZE 0.14 BY 0.16 ;
END MAS933

MACRO MAS934
   SIZE 0.14 BY 0.16 ;
END MAS934

MACRO MAS935
   SIZE 0.14 BY 0.16 ;
END MAS935

MACRO MAS936
   SIZE 0.14 BY 0.16 ;
END MAS936

MACRO MAS937
   SIZE 0.14 BY 0.16 ;
END MAS937

MACRO MAS938
   SIZE 0.14 BY 0.16 ;
END MAS938

MACRO MAS939
   SIZE 0.14 BY 0.16 ;
END MAS939

MACRO MAS940
   SIZE 0.14 BY 0.16 ;
END MAS940

MACRO MAS941
   SIZE 0.14 BY 0.16 ;
END MAS941

MACRO MAS942
   SIZE 0.14 BY 0.16 ;
END MAS942

MACRO MAS943
   SIZE 0.14 BY 0.16 ;
END MAS943

MACRO MAS944
   SIZE 0.14 BY 0.16 ;
END MAS944

MACRO MAS945
   SIZE 0.14 BY 0.16 ;
END MAS945

MACRO MAS946
   SIZE 0.14 BY 0.16 ;
END MAS946

MACRO MAS947
   SIZE 0.14 BY 0.16 ;
END MAS947

MACRO MAS948
   SIZE 0.14 BY 0.16 ;
END MAS948

MACRO MAS949
   SIZE 0.14 BY 0.16 ;
END MAS949

MACRO MAS950
   SIZE 0.14 BY 0.16 ;
END MAS950

MACRO MAS951
   SIZE 0.14 BY 0.16 ;
END MAS951

MACRO MAS952
   SIZE 0.14 BY 0.16 ;
END MAS952

MACRO MAS953
   SIZE 0.14 BY 0.16 ;
END MAS953

MACRO MAS954
   SIZE 0.14 BY 0.16 ;
END MAS954

MACRO MAS955
   SIZE 0.14 BY 0.16 ;
END MAS955

MACRO MAS956
   SIZE 0.14 BY 0.16 ;
END MAS956

MACRO MAS957
   SIZE 0.14 BY 0.16 ;
END MAS957

MACRO MAS958
   SIZE 0.14 BY 0.16 ;
END MAS958

MACRO MAS959
   SIZE 0.14 BY 0.16 ;
END MAS959

MACRO MAS960
   SIZE 0.14 BY 0.16 ;
END MAS960

MACRO MAS961
   SIZE 0.14 BY 0.16 ;
END MAS961

MACRO MAS962
   SIZE 0.14 BY 0.16 ;
END MAS962

MACRO MAS963
   SIZE 0.14 BY 0.16 ;
END MAS963

MACRO MAS964
   SIZE 0.14 BY 0.16 ;
END MAS964

MACRO MAS965
   SIZE 0.14 BY 0.16 ;
END MAS965

MACRO MAS966
   SIZE 0.14 BY 0.16 ;
END MAS966

MACRO MAS967
   SIZE 0.14 BY 0.16 ;
END MAS967

MACRO MAS968
   SIZE 0.14 BY 0.16 ;
END MAS968

MACRO MAS969
   SIZE 0.14 BY 0.16 ;
END MAS969

MACRO MAS970
   SIZE 0.14 BY 0.16 ;
END MAS970

MACRO MAS971
   SIZE 0.14 BY 0.16 ;
END MAS971

MACRO MAS972
   SIZE 0.14 BY 0.16 ;
END MAS972

MACRO MAS973
   SIZE 0.14 BY 0.16 ;
END MAS973

MACRO MAS974
   SIZE 0.14 BY 0.16 ;
END MAS974

MACRO MAS975
   SIZE 0.14 BY 0.16 ;
END MAS975

MACRO MAS976
   SIZE 0.14 BY 0.16 ;
END MAS976

MACRO MAS977
   SIZE 0.14 BY 0.16 ;
END MAS977

MACRO MAS978
   SIZE 0.14 BY 0.16 ;
END MAS978

MACRO MAS979
   SIZE 0.14 BY 0.16 ;
END MAS979

MACRO MAS980
   SIZE 0.14 BY 0.16 ;
END MAS980

MACRO MAS981
   SIZE 0.14 BY 0.16 ;
END MAS981

MACRO MAS982
   SIZE 0.14 BY 0.16 ;
END MAS982

MACRO MAS983
   SIZE 0.14 BY 0.16 ;
END MAS983

MACRO MAS984
   SIZE 0.14 BY 0.16 ;
END MAS984

MACRO MAS985
   SIZE 0.14 BY 0.16 ;
END MAS985

MACRO MAS986
   SIZE 0.14 BY 0.16 ;
END MAS986

MACRO MAS987
   SIZE 0.14 BY 0.16 ;
END MAS987

MACRO MAS988
   SIZE 0.14 BY 0.16 ;
END MAS988

MACRO MAS989
   SIZE 0.14 BY 0.16 ;
END MAS989

MACRO MAS990
   SIZE 0.14 BY 0.16 ;
END MAS990

MACRO MAS991
   SIZE 0.14 BY 0.16 ;
END MAS991

MACRO MAS992
   SIZE 0.14 BY 0.16 ;
END MAS992

MACRO MAS993
   SIZE 0.14 BY 0.16 ;
END MAS993

MACRO MAS994
   SIZE 0.14 BY 0.16 ;
END MAS994

MACRO MAS995
   SIZE 0.14 BY 0.16 ;
END MAS995

MACRO MAS996
   SIZE 0.14 BY 0.16 ;
END MAS996

MACRO MAS997
   SIZE 0.14 BY 0.16 ;
END MAS997

MACRO MAS998
   SIZE 0.14 BY 0.16 ;
END MAS998

MACRO MAS999
   SIZE 0.14 BY 0.16 ;
END MAS999

MACRO MAS1000
   SIZE 0.14 BY 0.16 ;
END MAS1000

MACRO MAS1001
   SIZE 0.14 BY 0.16 ;
END MAS1001

MACRO MAS1002
   SIZE 0.14 BY 0.16 ;
END MAS1002

MACRO MAS1003
   SIZE 0.14 BY 0.16 ;
END MAS1003

MACRO MAS1004
   SIZE 0.14 BY 0.16 ;
END MAS1004

MACRO MAS1005
   SIZE 0.14 BY 0.16 ;
END MAS1005

MACRO MAS1006
   SIZE 0.14 BY 0.16 ;
END MAS1006

MACRO MAS1007
   SIZE 0.14 BY 0.16 ;
END MAS1007

MACRO MAS1008
   SIZE 0.14 BY 0.16 ;
END MAS1008

MACRO MAS1009
   SIZE 0.14 BY 0.16 ;
END MAS1009

MACRO MAS1010
   SIZE 0.14 BY 0.16 ;
END MAS1010

MACRO MAS1011
   SIZE 0.14 BY 0.16 ;
END MAS1011

MACRO MAS1012
   SIZE 0.14 BY 0.16 ;
END MAS1012

MACRO MAS1013
   SIZE 0.14 BY 0.16 ;
END MAS1013

MACRO MAS1014
   SIZE 0.14 BY 0.16 ;
END MAS1014

MACRO MAS1015
   SIZE 0.14 BY 0.16 ;
END MAS1015

MACRO MAS1016
   SIZE 0.14 BY 0.16 ;
END MAS1016

MACRO MAS1017
   SIZE 0.14 BY 0.16 ;
END MAS1017

MACRO MAS1018
   SIZE 0.14 BY 0.16 ;
END MAS1018

MACRO MAS1019
   SIZE 0.14 BY 0.16 ;
END MAS1019

MACRO MAS1020
   SIZE 0.14 BY 0.16 ;
END MAS1020

MACRO MAS1021
   SIZE 0.14 BY 0.16 ;
END MAS1021

MACRO MAS1022
   SIZE 0.14 BY 0.16 ;
END MAS1022

MACRO MAS1023
   SIZE 0.14 BY 0.16 ;
END MAS1023

MACRO MAS1024
   SIZE 0.14 BY 0.16 ;
END MAS1024

MACRO MAS1025
   SIZE 0.14 BY 0.16 ;
END MAS1025

MACRO MAS1026
   SIZE 0.14 BY 0.16 ;
END MAS1026

MACRO MAS1027
   SIZE 0.14 BY 0.16 ;
END MAS1027

MACRO MAS1028
   SIZE 0.14 BY 0.16 ;
END MAS1028

MACRO MAS1029
   SIZE 0.14 BY 0.16 ;
END MAS1029

MACRO MAS1030
   SIZE 0.14 BY 0.16 ;
END MAS1030

MACRO MAS1031
   SIZE 0.14 BY 0.16 ;
END MAS1031

MACRO MAS1032
   SIZE 0.14 BY 0.16 ;
END MAS1032

MACRO MAS1033
   SIZE 0.14 BY 0.16 ;
END MAS1033

MACRO MAS1034
   SIZE 0.14 BY 0.16 ;
END MAS1034

MACRO MAS1035
   SIZE 0.14 BY 0.16 ;
END MAS1035

MACRO MAS1036
   SIZE 0.14 BY 0.16 ;
END MAS1036

MACRO MAS1037
   SIZE 0.14 BY 0.16 ;
END MAS1037

MACRO MAS1038
   SIZE 0.14 BY 0.16 ;
END MAS1038

MACRO MAS1039
   SIZE 0.14 BY 0.16 ;
END MAS1039

MACRO MAS1040
   SIZE 0.14 BY 0.16 ;
END MAS1040

MACRO MAS1041
   SIZE 0.14 BY 0.16 ;
END MAS1041

MACRO MAS1042
   SIZE 0.14 BY 0.16 ;
END MAS1042

MACRO MAS1043
   SIZE 0.14 BY 0.16 ;
END MAS1043

MACRO MAS1044
   SIZE 0.14 BY 0.16 ;
END MAS1044

MACRO MAS1045
   SIZE 0.14 BY 0.16 ;
END MAS1045

MACRO MAS1046
   SIZE 0.14 BY 0.16 ;
END MAS1046

MACRO MAS1047
   SIZE 0.14 BY 0.16 ;
END MAS1047

MACRO MAS1048
   SIZE 0.14 BY 0.16 ;
END MAS1048

MACRO MAS1049
   SIZE 0.14 BY 0.16 ;
END MAS1049

MACRO MAS1050
   SIZE 0.14 BY 0.16 ;
END MAS1050

MACRO MAS1051
   SIZE 0.14 BY 0.16 ;
END MAS1051

MACRO MAS1052
   SIZE 0.14 BY 0.16 ;
END MAS1052

MACRO MAS1053
   SIZE 0.14 BY 0.16 ;
END MAS1053

MACRO MAS1054
   SIZE 0.14 BY 0.16 ;
END MAS1054

MACRO MAS1055
   SIZE 0.14 BY 0.16 ;
END MAS1055

MACRO MAS1056
   SIZE 0.14 BY 0.16 ;
END MAS1056

MACRO MAS1057
   SIZE 0.14 BY 0.16 ;
END MAS1057

MACRO MAS1058
   SIZE 0.14 BY 0.16 ;
END MAS1058

MACRO MAS1059
   SIZE 0.14 BY 0.16 ;
END MAS1059

MACRO MAS1060
   SIZE 0.14 BY 0.16 ;
END MAS1060

MACRO MAS1061
   SIZE 0.14 BY 0.16 ;
END MAS1061

MACRO MAS1062
   SIZE 0.14 BY 0.16 ;
END MAS1062

MACRO MAS1063
   SIZE 0.14 BY 0.16 ;
END MAS1063

MACRO MAS1064
   SIZE 0.14 BY 0.16 ;
END MAS1064

MACRO MAS1065
   SIZE 0.14 BY 0.16 ;
END MAS1065

MACRO MAS1066
   SIZE 0.14 BY 0.16 ;
END MAS1066

MACRO MAS1067
   SIZE 0.14 BY 0.16 ;
END MAS1067

MACRO MAS1068
   SIZE 0.14 BY 0.16 ;
END MAS1068

MACRO MAS1069
   SIZE 0.14 BY 0.16 ;
END MAS1069

MACRO MAS1070
   SIZE 0.14 BY 0.16 ;
END MAS1070

MACRO MAS1071
   SIZE 0.14 BY 0.16 ;
END MAS1071

MACRO MAS1072
   SIZE 0.14 BY 0.16 ;
END MAS1072

MACRO MAS1073
   SIZE 0.14 BY 0.16 ;
END MAS1073

MACRO MAS1074
   SIZE 0.14 BY 0.16 ;
END MAS1074

MACRO MAS1075
   SIZE 0.14 BY 0.16 ;
END MAS1075

MACRO MAS1076
   SIZE 0.14 BY 0.16 ;
END MAS1076

MACRO MAS1077
   SIZE 0.14 BY 0.16 ;
END MAS1077

MACRO MAS1078
   SIZE 0.14 BY 0.16 ;
END MAS1078

MACRO MAS1079
   SIZE 0.14 BY 0.16 ;
END MAS1079

MACRO MAS1080
   SIZE 0.14 BY 0.16 ;
END MAS1080

MACRO MAS1081
   SIZE 0.14 BY 0.16 ;
END MAS1081

MACRO MAS1082
   SIZE 0.14 BY 0.16 ;
END MAS1082

MACRO MAS1083
   SIZE 0.14 BY 0.16 ;
END MAS1083

MACRO MAS1084
   SIZE 0.14 BY 0.16 ;
END MAS1084

MACRO MAS1085
   SIZE 0.14 BY 0.16 ;
END MAS1085

MACRO MAS1086
   SIZE 0.14 BY 0.16 ;
END MAS1086

MACRO MAS1087
   SIZE 0.14 BY 0.16 ;
END MAS1087

MACRO MAS1088
   SIZE 0.14 BY 0.16 ;
END MAS1088

MACRO MAS1089
   SIZE 0.14 BY 0.16 ;
END MAS1089

MACRO MAS1090
   SIZE 0.14 BY 0.16 ;
END MAS1090

MACRO MAS1091
   SIZE 0.14 BY 0.16 ;
END MAS1091

MACRO MAS1092
   SIZE 0.14 BY 0.16 ;
END MAS1092

MACRO MAS1093
   SIZE 0.14 BY 0.16 ;
END MAS1093

MACRO MAS1094
   SIZE 0.14 BY 0.16 ;
END MAS1094

MACRO MAS1095
   SIZE 0.14 BY 0.16 ;
END MAS1095

MACRO MAS1096
   SIZE 0.14 BY 0.16 ;
END MAS1096

MACRO MAS1097
   SIZE 0.14 BY 0.16 ;
END MAS1097

MACRO MAS1098
   SIZE 0.14 BY 0.16 ;
END MAS1098

MACRO MAS1099
   SIZE 0.14 BY 0.16 ;
END MAS1099

MACRO MAS1100
   SIZE 0.14 BY 0.16 ;
END MAS1100

MACRO MAS1101
   SIZE 0.14 BY 0.16 ;
END MAS1101

MACRO MAS1102
   SIZE 0.14 BY 0.16 ;
END MAS1102

MACRO MAS1103
   SIZE 0.14 BY 0.16 ;
END MAS1103

MACRO MAS1104
   SIZE 0.14 BY 0.16 ;
END MAS1104

MACRO MAS1105
   SIZE 0.14 BY 0.16 ;
END MAS1105

MACRO MAS1106
   SIZE 0.14 BY 0.16 ;
END MAS1106

MACRO MAS1107
   SIZE 0.14 BY 0.16 ;
END MAS1107

MACRO MAS1108
   SIZE 0.14 BY 0.16 ;
END MAS1108

MACRO MAS1109
   SIZE 0.14 BY 0.16 ;
END MAS1109

MACRO MAS1110
   SIZE 0.14 BY 0.16 ;
END MAS1110

MACRO MAS1111
   SIZE 0.14 BY 0.16 ;
END MAS1111

MACRO MAS1112
   SIZE 0.14 BY 0.16 ;
END MAS1112

MACRO MAS1113
   SIZE 0.14 BY 0.16 ;
END MAS1113

MACRO MAS1114
   SIZE 0.14 BY 0.16 ;
END MAS1114

MACRO MAS1115
   SIZE 0.14 BY 0.16 ;
END MAS1115

MACRO MAS1116
   SIZE 0.14 BY 0.16 ;
END MAS1116

MACRO MAS1117
   SIZE 0.14 BY 0.16 ;
END MAS1117

MACRO MAS1118
   SIZE 0.14 BY 0.16 ;
END MAS1118

MACRO MAS1119
   SIZE 0.14 BY 0.16 ;
END MAS1119

MACRO MAS1120
   SIZE 0.14 BY 0.16 ;
END MAS1120

MACRO MAS1121
   SIZE 0.14 BY 0.16 ;
END MAS1121

MACRO MAS1122
   SIZE 0.14 BY 0.16 ;
END MAS1122

MACRO MAS1123
   SIZE 0.14 BY 0.16 ;
END MAS1123

MACRO MAS1124
   SIZE 0.14 BY 0.16 ;
END MAS1124

MACRO MAS1125
   SIZE 0.14 BY 0.16 ;
END MAS1125

MACRO MAS1126
   SIZE 0.14 BY 0.16 ;
END MAS1126

MACRO MAS1127
   SIZE 0.14 BY 0.16 ;
END MAS1127

MACRO MAS1128
   SIZE 0.14 BY 0.16 ;
END MAS1128

MACRO MAS1129
   SIZE 0.14 BY 0.16 ;
END MAS1129

MACRO MAS1130
   SIZE 0.14 BY 0.16 ;
END MAS1130

MACRO MAS1131
   SIZE 0.14 BY 0.16 ;
END MAS1131

MACRO MAS1132
   SIZE 0.14 BY 0.16 ;
END MAS1132

MACRO MAS1133
   SIZE 0.14 BY 0.16 ;
END MAS1133

MACRO MAS1134
   SIZE 0.14 BY 0.16 ;
END MAS1134

MACRO MAS1135
   SIZE 0.14 BY 0.16 ;
END MAS1135

MACRO MAS1136
   SIZE 0.14 BY 0.16 ;
END MAS1136

MACRO MAS1137
   SIZE 0.14 BY 0.16 ;
END MAS1137

MACRO MAS1138
   SIZE 0.14 BY 0.16 ;
END MAS1138

MACRO MAS1139
   SIZE 0.14 BY 0.16 ;
END MAS1139

MACRO MAS1140
   SIZE 0.14 BY 0.16 ;
END MAS1140

MACRO MAS1141
   SIZE 0.14 BY 0.16 ;
END MAS1141

MACRO MAS1142
   SIZE 0.14 BY 0.16 ;
END MAS1142

MACRO MAS1143
   SIZE 0.14 BY 0.16 ;
END MAS1143

MACRO MAS1144
   SIZE 0.14 BY 0.16 ;
END MAS1144

MACRO MAS1145
   SIZE 0.14 BY 0.16 ;
END MAS1145

MACRO MAS1146
   SIZE 0.14 BY 0.16 ;
END MAS1146

MACRO MAS1147
   SIZE 0.14 BY 0.16 ;
END MAS1147

MACRO MAS1148
   SIZE 0.14 BY 0.16 ;
END MAS1148

MACRO MAS1149
   SIZE 0.14 BY 0.16 ;
END MAS1149

MACRO MAS1150
   SIZE 0.14 BY 0.16 ;
END MAS1150

MACRO MAS1151
   SIZE 0.14 BY 0.16 ;
END MAS1151

MACRO MAS1152
   SIZE 0.14 BY 0.16 ;
END MAS1152

MACRO MAS1153
   SIZE 0.14 BY 0.16 ;
END MAS1153

MACRO MAS1154
   SIZE 0.14 BY 0.16 ;
END MAS1154

MACRO MAS1155
   SIZE 0.14 BY 0.16 ;
END MAS1155

MACRO MAS1156
   SIZE 0.14 BY 0.16 ;
END MAS1156

MACRO MAS1157
   SIZE 0.14 BY 0.16 ;
END MAS1157

MACRO MAS1158
   SIZE 0.14 BY 0.16 ;
END MAS1158

MACRO MAS1159
   SIZE 0.14 BY 0.16 ;
END MAS1159

MACRO MAS1160
   SIZE 0.14 BY 0.16 ;
END MAS1160

MACRO MAS1161
   SIZE 0.14 BY 0.16 ;
END MAS1161

MACRO MAS1162
   SIZE 0.14 BY 0.16 ;
END MAS1162

MACRO MAS1163
   SIZE 0.14 BY 0.16 ;
END MAS1163

MACRO MAS1164
   SIZE 0.14 BY 0.16 ;
END MAS1164

MACRO MAS1165
   SIZE 0.14 BY 0.16 ;
END MAS1165

MACRO MAS1166
   SIZE 0.14 BY 0.16 ;
END MAS1166

MACRO MAS1167
   SIZE 0.14 BY 0.16 ;
END MAS1167

MACRO MAS1168
   SIZE 0.14 BY 0.16 ;
END MAS1168

MACRO MAS1169
   SIZE 0.14 BY 0.16 ;
END MAS1169

MACRO MAS1170
   SIZE 0.14 BY 0.16 ;
END MAS1170

MACRO MAS1171
   SIZE 0.14 BY 0.16 ;
END MAS1171

MACRO MAS1172
   SIZE 0.14 BY 0.16 ;
END MAS1172

MACRO MAS1173
   SIZE 0.14 BY 0.16 ;
END MAS1173

MACRO MAS1174
   SIZE 0.14 BY 0.16 ;
END MAS1174

MACRO MAS1175
   SIZE 0.14 BY 0.16 ;
END MAS1175

MACRO MAS1176
   SIZE 0.14 BY 0.16 ;
END MAS1176

MACRO MAS1177
   SIZE 0.14 BY 0.16 ;
END MAS1177

MACRO MAS1178
   SIZE 0.14 BY 0.16 ;
END MAS1178

MACRO MAS1179
   SIZE 0.14 BY 0.16 ;
END MAS1179

MACRO MAS1180
   SIZE 0.14 BY 0.16 ;
END MAS1180

MACRO MAS1181
   SIZE 0.14 BY 0.16 ;
END MAS1181

MACRO MAS1182
   SIZE 0.14 BY 0.16 ;
END MAS1182

MACRO MAS1183
   SIZE 0.14 BY 0.16 ;
END MAS1183

MACRO MAS1184
   SIZE 0.14 BY 0.16 ;
END MAS1184

MACRO MAS1185
   SIZE 0.14 BY 0.16 ;
END MAS1185

MACRO MAS1186
   SIZE 0.14 BY 0.16 ;
END MAS1186

MACRO MAS1187
   SIZE 0.14 BY 0.16 ;
END MAS1187

MACRO MAS1188
   SIZE 0.14 BY 0.16 ;
END MAS1188

MACRO MAS1189
   SIZE 0.14 BY 0.16 ;
END MAS1189

MACRO MAS1190
   SIZE 0.14 BY 0.16 ;
END MAS1190

MACRO MAS1191
   SIZE 0.14 BY 0.16 ;
END MAS1191

MACRO MAS1192
   SIZE 0.14 BY 0.16 ;
END MAS1192

MACRO MAS1193
   SIZE 0.14 BY 0.16 ;
END MAS1193

MACRO MAS1194
   SIZE 0.14 BY 0.16 ;
END MAS1194

MACRO MAS1195
   SIZE 0.14 BY 0.16 ;
END MAS1195

MACRO MAS1196
   SIZE 0.14 BY 0.16 ;
END MAS1196

MACRO MAS1197
   SIZE 0.14 BY 0.16 ;
END MAS1197

MACRO MAS1198
   SIZE 0.14 BY 0.16 ;
END MAS1198

MACRO MAS1199
   SIZE 0.14 BY 0.16 ;
END MAS1199

MACRO MAS1200
   SIZE 0.14 BY 0.16 ;
END MAS1200

MACRO MAS1201
   SIZE 0.14 BY 0.16 ;
END MAS1201

MACRO MAS1202
   SIZE 0.14 BY 0.16 ;
END MAS1202

MACRO MAS1203
   SIZE 0.14 BY 0.16 ;
END MAS1203

MACRO MAS1204
   SIZE 0.14 BY 0.16 ;
END MAS1204

MACRO MAS1205
   SIZE 0.14 BY 0.16 ;
END MAS1205

MACRO MAS1206
   SIZE 0.14 BY 0.16 ;
END MAS1206

MACRO MAS1207
   SIZE 0.14 BY 0.16 ;
END MAS1207

MACRO MAS1208
   SIZE 0.14 BY 0.16 ;
END MAS1208

MACRO MAS1209
   SIZE 0.14 BY 0.16 ;
END MAS1209

MACRO MAS1210
   SIZE 0.14 BY 0.16 ;
END MAS1210

MACRO MAS1211
   SIZE 0.14 BY 0.16 ;
END MAS1211

MACRO MAS1212
   SIZE 0.14 BY 0.16 ;
END MAS1212

MACRO MAS1213
   SIZE 0.14 BY 0.16 ;
END MAS1213

MACRO MAS1214
   SIZE 0.14 BY 0.16 ;
END MAS1214

MACRO MAS1215
   SIZE 0.14 BY 0.16 ;
END MAS1215

MACRO MAS1216
   SIZE 0.14 BY 0.16 ;
END MAS1216

MACRO MAS1217
   SIZE 0.14 BY 0.16 ;
END MAS1217

MACRO MAS1218
   SIZE 0.14 BY 0.16 ;
END MAS1218

MACRO MAS1219
   SIZE 0.14 BY 0.16 ;
END MAS1219

MACRO MAS1220
   SIZE 0.14 BY 0.16 ;
END MAS1220

MACRO MAS1221
   SIZE 0.14 BY 0.16 ;
END MAS1221

MACRO MAS1222
   SIZE 0.14 BY 0.16 ;
END MAS1222

MACRO MAS1223
   SIZE 0.14 BY 0.16 ;
END MAS1223

MACRO MAS1224
   SIZE 0.14 BY 0.16 ;
END MAS1224

MACRO MAS1225
   SIZE 0.14 BY 0.16 ;
END MAS1225

MACRO MAS1226
   SIZE 0.14 BY 0.16 ;
END MAS1226

MACRO MAS1227
   SIZE 0.14 BY 0.16 ;
END MAS1227

MACRO MAS1228
   SIZE 0.14 BY 0.16 ;
END MAS1228

MACRO MAS1229
   SIZE 0.14 BY 0.16 ;
END MAS1229

MACRO MAS1230
   SIZE 0.14 BY 0.16 ;
END MAS1230

MACRO MAS1231
   SIZE 0.14 BY 0.16 ;
END MAS1231

MACRO MAS1232
   SIZE 0.14 BY 0.16 ;
END MAS1232

MACRO MAS1233
   SIZE 0.14 BY 0.16 ;
END MAS1233

MACRO MAS1234
   SIZE 0.14 BY 0.16 ;
END MAS1234

MACRO MAS1235
   SIZE 0.14 BY 0.16 ;
END MAS1235

MACRO MAS1236
   SIZE 0.14 BY 0.16 ;
END MAS1236

MACRO MAS1237
   SIZE 0.14 BY 0.16 ;
END MAS1237

MACRO MAS1238
   SIZE 0.14 BY 0.16 ;
END MAS1238

MACRO MAS1239
   SIZE 0.14 BY 0.16 ;
END MAS1239

MACRO MAS1240
   SIZE 0.14 BY 0.16 ;
END MAS1240

MACRO MAS1241
   SIZE 0.14 BY 0.16 ;
END MAS1241

MACRO MAS1242
   SIZE 0.14 BY 0.16 ;
END MAS1242

MACRO MAS1243
   SIZE 0.14 BY 0.16 ;
END MAS1243

MACRO MAS1244
   SIZE 0.14 BY 0.16 ;
END MAS1244

MACRO MAS1245
   SIZE 0.14 BY 0.16 ;
END MAS1245

MACRO MAS1246
   SIZE 0.14 BY 0.16 ;
END MAS1246

MACRO MAS1247
   SIZE 0.14 BY 0.16 ;
END MAS1247

MACRO MAS1248
   SIZE 0.14 BY 0.16 ;
END MAS1248

MACRO MAS1249
   SIZE 0.14 BY 0.16 ;
END MAS1249

MACRO MAS1250
   SIZE 0.14 BY 0.16 ;
END MAS1250

MACRO MAS1251
   SIZE 0.14 BY 0.16 ;
END MAS1251

MACRO MAS1252
   SIZE 0.14 BY 0.16 ;
END MAS1252

MACRO MAS1253
   SIZE 0.14 BY 0.16 ;
END MAS1253

MACRO MAS1254
   SIZE 0.14 BY 0.16 ;
END MAS1254

MACRO MAS1255
   SIZE 0.14 BY 0.16 ;
END MAS1255

MACRO MAS1256
   SIZE 0.14 BY 0.16 ;
END MAS1256

MACRO MAS1257
   SIZE 0.14 BY 0.16 ;
END MAS1257

MACRO MAS1258
   SIZE 0.14 BY 0.16 ;
END MAS1258

MACRO MAS1259
   SIZE 0.14 BY 0.16 ;
END MAS1259

MACRO MAS1260
   SIZE 0.14 BY 0.16 ;
END MAS1260

MACRO MAS1261
   SIZE 0.14 BY 0.16 ;
END MAS1261

MACRO MAS1262
   SIZE 0.14 BY 0.16 ;
END MAS1262

MACRO MAS1263
   SIZE 0.14 BY 0.16 ;
END MAS1263

MACRO MAS1264
   SIZE 0.14 BY 0.16 ;
END MAS1264

MACRO MAS1265
   SIZE 0.14 BY 0.16 ;
END MAS1265

MACRO MAS1266
   SIZE 0.14 BY 0.16 ;
END MAS1266

MACRO MAS1267
   SIZE 0.14 BY 0.16 ;
END MAS1267

MACRO MAS1268
   SIZE 0.14 BY 0.16 ;
END MAS1268

MACRO MAS1269
   SIZE 0.14 BY 0.16 ;
END MAS1269

MACRO MAS1270
   SIZE 0.14 BY 0.16 ;
END MAS1270

MACRO MAS1271
   SIZE 0.14 BY 0.16 ;
END MAS1271

MACRO MAS1272
   SIZE 0.14 BY 0.16 ;
END MAS1272

MACRO MAS1273
   SIZE 0.14 BY 0.16 ;
END MAS1273

MACRO MAS1274
   SIZE 0.14 BY 0.16 ;
END MAS1274

MACRO MAS1275
   SIZE 0.14 BY 0.16 ;
END MAS1275

MACRO MAS1276
   SIZE 0.14 BY 0.16 ;
END MAS1276

MACRO MAS1277
   SIZE 0.14 BY 0.16 ;
END MAS1277

MACRO MAS1278
   SIZE 0.14 BY 0.16 ;
END MAS1278

MACRO MAS1279
   SIZE 0.14 BY 0.16 ;
END MAS1279

MACRO MAS1280
   SIZE 0.14 BY 0.16 ;
END MAS1280

MACRO MAS1281
   SIZE 0.14 BY 0.16 ;
END MAS1281

MACRO MAS1282
   SIZE 0.14 BY 0.16 ;
END MAS1282

MACRO MAS1283
   SIZE 0.14 BY 0.16 ;
END MAS1283

MACRO MAS1284
   SIZE 0.14 BY 0.16 ;
END MAS1284

MACRO MAS1285
   SIZE 0.14 BY 0.16 ;
END MAS1285

MACRO MAS1286
   SIZE 0.14 BY 0.16 ;
END MAS1286

MACRO MAS1287
   SIZE 0.14 BY 0.16 ;
END MAS1287

MACRO MAS1288
   SIZE 0.14 BY 0.16 ;
END MAS1288

MACRO MAS1289
   SIZE 0.14 BY 0.16 ;
END MAS1289

MACRO MAS1290
   SIZE 0.14 BY 0.16 ;
END MAS1290

MACRO MAS1291
   SIZE 0.14 BY 0.16 ;
END MAS1291

MACRO MAS1292
   SIZE 0.14 BY 0.16 ;
END MAS1292

MACRO MAS1293
   SIZE 0.14 BY 0.16 ;
END MAS1293

MACRO MAS1294
   SIZE 0.14 BY 0.16 ;
END MAS1294

MACRO MAS1295
   SIZE 0.14 BY 0.16 ;
END MAS1295

MACRO MAS1296
   SIZE 0.14 BY 0.16 ;
END MAS1296

MACRO MAS1297
   SIZE 0.14 BY 0.16 ;
END MAS1297

MACRO MAS1298
   SIZE 0.14 BY 0.16 ;
END MAS1298

MACRO MAS1299
   SIZE 0.14 BY 0.16 ;
END MAS1299

MACRO MAS1300
   SIZE 0.14 BY 0.16 ;
END MAS1300

MACRO MAS1301
   SIZE 0.14 BY 0.16 ;
END MAS1301

MACRO MAS1302
   SIZE 0.14 BY 0.16 ;
END MAS1302

MACRO MAS1303
   SIZE 0.14 BY 0.16 ;
END MAS1303

MACRO MAS1304
   SIZE 0.14 BY 0.16 ;
END MAS1304

MACRO MAS1305
   SIZE 0.14 BY 0.16 ;
END MAS1305

MACRO MAS1306
   SIZE 0.14 BY 0.16 ;
END MAS1306

MACRO MAS1307
   SIZE 0.14 BY 0.16 ;
END MAS1307

MACRO MAS1308
   SIZE 0.14 BY 0.16 ;
END MAS1308

MACRO MAS1309
   SIZE 0.14 BY 0.16 ;
END MAS1309

MACRO MAS1310
   SIZE 0.14 BY 0.16 ;
END MAS1310

MACRO MAS1311
   SIZE 0.14 BY 0.16 ;
END MAS1311

MACRO MAS1312
   SIZE 0.14 BY 0.16 ;
END MAS1312

MACRO MAS1313
   SIZE 0.14 BY 0.16 ;
END MAS1313

MACRO MAS1314
   SIZE 0.14 BY 0.16 ;
END MAS1314

MACRO MAS1315
   SIZE 0.14 BY 0.16 ;
END MAS1315

MACRO MAS1316
   SIZE 0.14 BY 0.16 ;
END MAS1316

MACRO MAS1317
   SIZE 0.14 BY 0.16 ;
END MAS1317

MACRO MAS1318
   SIZE 0.14 BY 0.16 ;
END MAS1318

MACRO MAS1319
   SIZE 0.14 BY 0.16 ;
END MAS1319

MACRO MAS1320
   SIZE 0.14 BY 0.16 ;
END MAS1320

MACRO MAS1321
   SIZE 0.14 BY 0.16 ;
END MAS1321

MACRO MAS1322
   SIZE 0.14 BY 0.16 ;
END MAS1322

MACRO MAS1323
   SIZE 0.14 BY 0.16 ;
END MAS1323

MACRO MAS1324
   SIZE 0.14 BY 0.16 ;
END MAS1324

MACRO MAS1325
   SIZE 0.14 BY 0.16 ;
END MAS1325

MACRO MAS1326
   SIZE 0.14 BY 0.16 ;
END MAS1326

MACRO MAS1327
   SIZE 0.14 BY 0.16 ;
END MAS1327

MACRO MAS1328
   SIZE 0.14 BY 0.16 ;
END MAS1328

MACRO MAS1329
   SIZE 0.14 BY 0.16 ;
END MAS1329

MACRO MAS1330
   SIZE 0.14 BY 0.16 ;
END MAS1330

MACRO MAS1331
   SIZE 0.14 BY 0.16 ;
END MAS1331

MACRO MAS1332
   SIZE 0.14 BY 0.16 ;
END MAS1332

MACRO MAS1333
   SIZE 0.14 BY 0.16 ;
END MAS1333

MACRO MAS1334
   SIZE 0.14 BY 0.16 ;
END MAS1334

MACRO MAS1335
   SIZE 0.14 BY 0.16 ;
END MAS1335

MACRO MAS1336
   SIZE 0.14 BY 0.16 ;
END MAS1336

MACRO MAS1337
   SIZE 0.14 BY 0.16 ;
END MAS1337

MACRO MAS1338
   SIZE 0.14 BY 0.16 ;
END MAS1338

MACRO MAS1339
   SIZE 0.14 BY 0.16 ;
END MAS1339

MACRO MAS1340
   SIZE 0.14 BY 0.16 ;
END MAS1340

MACRO MAS1341
   SIZE 0.14 BY 0.16 ;
END MAS1341

MACRO MAS1342
   SIZE 0.14 BY 0.16 ;
END MAS1342

MACRO MAS1343
   SIZE 0.14 BY 0.16 ;
END MAS1343

MACRO MAS1344
   SIZE 0.14 BY 0.16 ;
END MAS1344

MACRO MAS1345
   SIZE 0.14 BY 0.16 ;
END MAS1345

MACRO MAS1346
   SIZE 0.14 BY 0.16 ;
END MAS1346

MACRO MAS1347
   SIZE 0.14 BY 0.16 ;
END MAS1347

MACRO MAS1348
   SIZE 0.14 BY 0.16 ;
END MAS1348

MACRO MAS1349
   SIZE 0.14 BY 0.16 ;
END MAS1349

MACRO MAS1350
   SIZE 0.14 BY 0.16 ;
END MAS1350

MACRO MAS1351
   SIZE 0.14 BY 0.16 ;
END MAS1351

MACRO MAS1352
   SIZE 0.14 BY 0.16 ;
END MAS1352

MACRO MAS1353
   SIZE 0.14 BY 0.16 ;
END MAS1353

MACRO MAS1354
   SIZE 0.14 BY 0.16 ;
END MAS1354

MACRO MAS1355
   SIZE 0.14 BY 0.16 ;
END MAS1355

MACRO MAS1356
   SIZE 0.14 BY 0.16 ;
END MAS1356

MACRO MAS1357
   SIZE 0.14 BY 0.16 ;
END MAS1357

MACRO MAS1358
   SIZE 0.14 BY 0.16 ;
END MAS1358

MACRO MAS1359
   SIZE 0.14 BY 0.16 ;
END MAS1359

MACRO MAS1360
   SIZE 0.14 BY 0.16 ;
END MAS1360

MACRO MAS1361
   SIZE 0.14 BY 0.16 ;
END MAS1361

MACRO MAS1362
   SIZE 0.14 BY 0.16 ;
END MAS1362

MACRO MAS1363
   SIZE 0.14 BY 0.16 ;
END MAS1363

MACRO MAS1364
   SIZE 0.14 BY 0.16 ;
END MAS1364

MACRO MAS1365
   SIZE 0.14 BY 0.16 ;
END MAS1365

MACRO MAS1366
   SIZE 0.14 BY 0.16 ;
END MAS1366

MACRO MAS1367
   SIZE 0.14 BY 0.16 ;
END MAS1367

MACRO MAS1368
   SIZE 0.14 BY 0.16 ;
END MAS1368

MACRO MAS1369
   SIZE 0.14 BY 0.16 ;
END MAS1369

MACRO MAS1370
   SIZE 0.14 BY 0.16 ;
END MAS1370

MACRO MAS1371
   SIZE 0.14 BY 0.16 ;
END MAS1371

MACRO MAS1372
   SIZE 0.14 BY 0.16 ;
END MAS1372

MACRO MAS1373
   SIZE 0.14 BY 0.16 ;
END MAS1373

MACRO MAS1374
   SIZE 0.14 BY 0.16 ;
END MAS1374

MACRO MAS1375
   SIZE 0.14 BY 0.16 ;
END MAS1375

MACRO MAS1376
   SIZE 0.14 BY 0.16 ;
END MAS1376

MACRO MAS1377
   SIZE 0.14 BY 0.16 ;
END MAS1377

MACRO MAS1378
   SIZE 0.14 BY 0.16 ;
END MAS1378

MACRO MAS1379
   SIZE 0.14 BY 0.16 ;
END MAS1379

MACRO MAS1380
   SIZE 0.14 BY 0.16 ;
END MAS1380

MACRO MAS1381
   SIZE 0.14 BY 0.16 ;
END MAS1381

MACRO MAS1382
   SIZE 0.14 BY 0.16 ;
END MAS1382

MACRO MAS1383
   SIZE 0.14 BY 0.16 ;
END MAS1383

MACRO MAS1384
   SIZE 0.14 BY 0.16 ;
END MAS1384

MACRO MAS1385
   SIZE 0.14 BY 0.16 ;
END MAS1385

MACRO MAS1386
   SIZE 0.14 BY 0.16 ;
END MAS1386

MACRO MAS1387
   SIZE 0.14 BY 0.16 ;
END MAS1387

MACRO MAS1388
   SIZE 0.14 BY 0.16 ;
END MAS1388

MACRO MAS1389
   SIZE 0.14 BY 0.16 ;
END MAS1389

MACRO MAS1390
   SIZE 0.16 BY 0.16 ;
END MAS1390

MACRO MAS1391
   SIZE 0.16 BY 0.16 ;
END MAS1391

MACRO MAS1392
   SIZE 0.16 BY 0.16 ;
END MAS1392

MACRO MAS1393
   SIZE 0.16 BY 0.16 ;
END MAS1393

MACRO MAS1394
   SIZE 0.16 BY 0.16 ;
END MAS1394

MACRO MAS1395
   SIZE 0.16 BY 0.16 ;
END MAS1395

MACRO MAS1396
   SIZE 0.16 BY 0.16 ;
END MAS1396

MACRO MAS1397
   SIZE 0.16 BY 0.16 ;
END MAS1397

MACRO MAS1398
   SIZE 0.16 BY 0.16 ;
END MAS1398

MACRO MAS1399
   SIZE 0.16 BY 0.16 ;
END MAS1399

MACRO MAS1400
   SIZE 0.16 BY 0.16 ;
END MAS1400

MACRO MAS1401
   SIZE 0.16 BY 0.16 ;
END MAS1401

MACRO MAS1402
   SIZE 0.16 BY 0.16 ;
END MAS1402

MACRO MAS1403
   SIZE 0.16 BY 0.16 ;
END MAS1403

MACRO MAS1404
   SIZE 0.16 BY 0.16 ;
END MAS1404

MACRO MAS1405
   SIZE 0.16 BY 0.16 ;
END MAS1405

MACRO MAS1406
   SIZE 0.16 BY 0.16 ;
END MAS1406

MACRO MAS1407
   SIZE 0.16 BY 0.16 ;
END MAS1407

MACRO MAS1408
   SIZE 0.16 BY 0.16 ;
END MAS1408

MACRO MAS1409
   SIZE 0.16 BY 0.16 ;
END MAS1409

MACRO MAS1410
   SIZE 0.16 BY 0.16 ;
END MAS1410

MACRO MAS1411
   SIZE 0.16 BY 0.16 ;
END MAS1411

MACRO MAS1412
   SIZE 0.16 BY 0.16 ;
END MAS1412

MACRO MAS1413
   SIZE 0.16 BY 0.16 ;
END MAS1413

MACRO MAS1414
   SIZE 0.16 BY 0.16 ;
END MAS1414

MACRO MAS1415
   SIZE 0.16 BY 0.16 ;
END MAS1415

MACRO MAS1416
   SIZE 0.16 BY 0.16 ;
END MAS1416

MACRO MAS1417
   SIZE 0.16 BY 0.16 ;
END MAS1417

MACRO MAS1418
   SIZE 0.16 BY 0.16 ;
END MAS1418

MACRO MAS1419
   SIZE 0.16 BY 0.16 ;
END MAS1419

MACRO MAS1420
   SIZE 0.16 BY 0.16 ;
END MAS1420

MACRO MAS1421
   SIZE 0.16 BY 0.16 ;
END MAS1421

MACRO MAS1422
   SIZE 0.16 BY 0.16 ;
END MAS1422

MACRO MAS1423
   SIZE 0.16 BY 0.16 ;
END MAS1423

MACRO MAS1424
   SIZE 0.16 BY 0.16 ;
END MAS1424

MACRO MAS1425
   SIZE 0.16 BY 0.16 ;
END MAS1425

MACRO MAS1426
   SIZE 0.16 BY 0.16 ;
END MAS1426

MACRO MAS1427
   SIZE 0.16 BY 0.16 ;
END MAS1427

MACRO MAS1428
   SIZE 0.16 BY 0.16 ;
END MAS1428

MACRO MAS1429
   SIZE 0.16 BY 0.16 ;
END MAS1429

MACRO MAS1430
   SIZE 0.16 BY 0.16 ;
END MAS1430

MACRO MAS1431
   SIZE 0.16 BY 0.16 ;
END MAS1431

MACRO MAS1432
   SIZE 0.16 BY 0.16 ;
END MAS1432

MACRO MAS1433
   SIZE 0.16 BY 0.16 ;
END MAS1433

MACRO MAS1434
   SIZE 0.16 BY 0.16 ;
END MAS1434

MACRO MAS1435
   SIZE 0.16 BY 0.16 ;
END MAS1435

MACRO MAS1436
   SIZE 0.16 BY 0.16 ;
END MAS1436

MACRO MAS1437
   SIZE 0.16 BY 0.16 ;
END MAS1437

MACRO MAS1438
   SIZE 0.16 BY 0.16 ;
END MAS1438

MACRO MAS1439
   SIZE 0.16 BY 0.16 ;
END MAS1439

MACRO MAS1440
   SIZE 0.16 BY 0.16 ;
END MAS1440

MACRO MAS1441
   SIZE 0.16 BY 0.16 ;
END MAS1441

MACRO MAS1442
   SIZE 0.16 BY 0.16 ;
END MAS1442

MACRO MAS1443
   SIZE 0.16 BY 0.16 ;
END MAS1443

MACRO MAS1444
   SIZE 0.16 BY 0.16 ;
END MAS1444

MACRO MAS1445
   SIZE 0.16 BY 0.16 ;
END MAS1445

MACRO MAS1446
   SIZE 0.16 BY 0.16 ;
END MAS1446

MACRO MAS1447
   SIZE 0.16 BY 0.16 ;
END MAS1447

MACRO MAS1448
   SIZE 0.16 BY 0.16 ;
END MAS1448

MACRO MAS1449
   SIZE 0.16 BY 0.16 ;
END MAS1449

MACRO MAS1450
   SIZE 0.16 BY 0.16 ;
END MAS1450

MACRO MAS1451
   SIZE 0.16 BY 0.16 ;
END MAS1451

MACRO MAS1452
   SIZE 0.16 BY 0.16 ;
END MAS1452

MACRO MAS1453
   SIZE 0.16 BY 0.16 ;
END MAS1453

MACRO MAS1454
   SIZE 0.16 BY 0.16 ;
END MAS1454

MACRO MAS1455
   SIZE 0.16 BY 0.16 ;
END MAS1455

MACRO MAS1456
   SIZE 0.16 BY 0.16 ;
END MAS1456

MACRO MAS1457
   SIZE 0.16 BY 0.16 ;
END MAS1457

MACRO MAS1458
   SIZE 0.16 BY 0.16 ;
END MAS1458

MACRO MAS1459
   SIZE 0.16 BY 0.16 ;
END MAS1459

MACRO MAS1460
   SIZE 0.16 BY 0.16 ;
END MAS1460

MACRO MAS1461
   SIZE 0.16 BY 0.16 ;
END MAS1461

MACRO MAS1462
   SIZE 0.16 BY 0.16 ;
END MAS1462

MACRO MAS1463
   SIZE 0.16 BY 0.16 ;
END MAS1463

MACRO MAS1464
   SIZE 0.16 BY 0.16 ;
END MAS1464

MACRO MAS1465
   SIZE 0.16 BY 0.16 ;
END MAS1465

MACRO MAS1466
   SIZE 0.16 BY 0.16 ;
END MAS1466

MACRO MAS1467
   SIZE 0.16 BY 0.16 ;
END MAS1467

MACRO MAS1468
   SIZE 0.16 BY 0.16 ;
END MAS1468

MACRO MAS1469
   SIZE 0.16 BY 0.16 ;
END MAS1469

MACRO MAS1470
   SIZE 0.16 BY 0.16 ;
END MAS1470

MACRO MAS1471
   SIZE 0.16 BY 0.16 ;
END MAS1471

MACRO MAS1472
   SIZE 0.16 BY 0.16 ;
END MAS1472

MACRO MAS1473
   SIZE 0.16 BY 0.16 ;
END MAS1473

MACRO MAS1474
   SIZE 0.16 BY 0.16 ;
END MAS1474

MACRO MAS1475
   SIZE 0.16 BY 0.16 ;
END MAS1475

MACRO MAS1476
   SIZE 0.16 BY 0.16 ;
END MAS1476

MACRO MAS1477
   SIZE 0.16 BY 0.16 ;
END MAS1477

MACRO MAS1478
   SIZE 0.16 BY 0.16 ;
END MAS1478

MACRO MAS1479
   SIZE 0.16 BY 0.16 ;
END MAS1479

MACRO MAS1480
   SIZE 0.16 BY 0.16 ;
END MAS1480

MACRO MAS1481
   SIZE 0.16 BY 0.16 ;
END MAS1481

MACRO MAS1482
   SIZE 0.16 BY 0.16 ;
END MAS1482

MACRO MAS1483
   SIZE 0.16 BY 0.16 ;
END MAS1483

MACRO MAS1484
   SIZE 0.16 BY 0.16 ;
END MAS1484

MACRO MAS1485
   SIZE 0.16 BY 0.16 ;
END MAS1485

MACRO MAS1486
   SIZE 0.16 BY 0.16 ;
END MAS1486

MACRO MAS1487
   SIZE 0.16 BY 0.16 ;
END MAS1487

MACRO MAS1488
   SIZE 0.16 BY 0.16 ;
END MAS1488

MACRO MAS1489
   SIZE 0.16 BY 0.16 ;
END MAS1489

MACRO MAS1490
   SIZE 0.16 BY 0.16 ;
END MAS1490

MACRO MAS1491
   SIZE 0.16 BY 0.16 ;
END MAS1491

MACRO MAS1492
   SIZE 0.16 BY 0.16 ;
END MAS1492

MACRO MAS1493
   SIZE 0.16 BY 0.16 ;
END MAS1493

MACRO MAS1494
   SIZE 0.16 BY 0.16 ;
END MAS1494

MACRO MAS1495
   SIZE 0.16 BY 0.16 ;
END MAS1495

MACRO MAS1496
   SIZE 0.16 BY 0.16 ;
END MAS1496

MACRO MAS1497
   SIZE 0.16 BY 0.16 ;
END MAS1497

MACRO MAS1498
   SIZE 0.16 BY 0.16 ;
END MAS1498

MACRO MAS1499
   SIZE 0.16 BY 0.16 ;
END MAS1499

MACRO MAS1500
   SIZE 0.16 BY 0.16 ;
END MAS1500

MACRO MAS1501
   SIZE 0.16 BY 0.16 ;
END MAS1501

MACRO MAS1502
   SIZE 0.16 BY 0.16 ;
END MAS1502

MACRO MAS1503
   SIZE 0.16 BY 0.16 ;
END MAS1503

MACRO MAS1504
   SIZE 0.16 BY 0.16 ;
END MAS1504

MACRO MAS1505
   SIZE 0.16 BY 0.16 ;
END MAS1505

MACRO MAS1506
   SIZE 0.16 BY 0.16 ;
END MAS1506

MACRO MAS1507
   SIZE 0.16 BY 0.16 ;
END MAS1507

MACRO MAS1508
   SIZE 0.16 BY 0.16 ;
END MAS1508

MACRO MAS1509
   SIZE 0.16 BY 0.16 ;
END MAS1509

MACRO MAS1510
   SIZE 0.16 BY 0.16 ;
END MAS1510

MACRO MAS1511
   SIZE 0.16 BY 0.16 ;
END MAS1511

MACRO MAS1512
   SIZE 0.16 BY 0.16 ;
END MAS1512

MACRO MAS1513
   SIZE 0.16 BY 0.16 ;
END MAS1513

MACRO MAS1514
   SIZE 0.16 BY 0.16 ;
END MAS1514

MACRO MAS1515
   SIZE 0.16 BY 0.16 ;
END MAS1515

MACRO MAS1516
   SIZE 0.16 BY 0.16 ;
END MAS1516

MACRO MAS1517
   SIZE 0.16 BY 0.16 ;
END MAS1517

MACRO MAS1518
   SIZE 0.16 BY 0.16 ;
END MAS1518

MACRO MAS1519
   SIZE 0.16 BY 0.16 ;
END MAS1519

MACRO MAS1520
   SIZE 0.16 BY 0.16 ;
END MAS1520

MACRO MAS1521
   SIZE 0.16 BY 0.16 ;
END MAS1521

MACRO MAS1522
   SIZE 0.16 BY 0.16 ;
END MAS1522

MACRO MAS1523
   SIZE 0.16 BY 0.16 ;
END MAS1523

MACRO MAS1524
   SIZE 0.16 BY 0.16 ;
END MAS1524

MACRO MAS1525
   SIZE 0.16 BY 0.16 ;
END MAS1525

MACRO MAS1526
   SIZE 0.16 BY 0.16 ;
END MAS1526

MACRO MAS1527
   SIZE 0.16 BY 0.16 ;
END MAS1527

MACRO MAS1528
   SIZE 0.16 BY 0.16 ;
END MAS1528

MACRO MAS1529
   SIZE 0.16 BY 0.16 ;
END MAS1529

MACRO MAS1530
   SIZE 0.16 BY 0.16 ;
END MAS1530

MACRO MAS1531
   SIZE 0.16 BY 0.16 ;
END MAS1531

MACRO MAS1532
   SIZE 0.16 BY 0.16 ;
END MAS1532

MACRO MAS1533
   SIZE 0.16 BY 0.16 ;
END MAS1533

MACRO MAS1534
   SIZE 0.16 BY 0.16 ;
END MAS1534

MACRO MAS1535
   SIZE 0.16 BY 0.16 ;
END MAS1535

MACRO MAS1536
   SIZE 0.16 BY 0.16 ;
END MAS1536

MACRO MAS1537
   SIZE 0.16 BY 0.16 ;
END MAS1537

MACRO MAS1538
   SIZE 0.16 BY 0.16 ;
END MAS1538

MACRO MAS1539
   SIZE 0.16 BY 0.16 ;
END MAS1539

MACRO MAS1540
   SIZE 0.16 BY 0.16 ;
END MAS1540

MACRO MAS1541
   SIZE 0.16 BY 0.16 ;
END MAS1541

MACRO MAS1542
   SIZE 0.16 BY 0.16 ;
END MAS1542

MACRO MAS1543
   SIZE 0.16 BY 0.16 ;
END MAS1543

MACRO MAS1544
   SIZE 0.16 BY 0.16 ;
END MAS1544

MACRO MAS1545
   SIZE 0.16 BY 0.16 ;
END MAS1545

MACRO MAS1546
   SIZE 0.16 BY 0.16 ;
END MAS1546

MACRO MAS1547
   SIZE 0.16 BY 0.16 ;
END MAS1547

MACRO MAS1548
   SIZE 0.16 BY 0.16 ;
END MAS1548

MACRO MAS1549
   SIZE 0.16 BY 0.16 ;
END MAS1549

MACRO MAS1550
   SIZE 0.16 BY 0.16 ;
END MAS1550

MACRO MAS1551
   SIZE 0.16 BY 0.16 ;
END MAS1551

MACRO MAS1552
   SIZE 0.16 BY 0.16 ;
END MAS1552

MACRO MAS1553
   SIZE 0.16 BY 0.16 ;
END MAS1553

MACRO MAS1554
   SIZE 0.16 BY 0.16 ;
END MAS1554

MACRO MAS1555
   SIZE 0.16 BY 0.16 ;
END MAS1555

MACRO MAS1556
   SIZE 0.16 BY 0.16 ;
END MAS1556

MACRO MAS1557
   SIZE 0.16 BY 0.16 ;
END MAS1557

MACRO MAS1558
   SIZE 0.16 BY 0.16 ;
END MAS1558

MACRO MAS1559
   SIZE 0.16 BY 0.16 ;
END MAS1559

MACRO MAS1560
   SIZE 0.16 BY 0.16 ;
END MAS1560

MACRO MAS1561
   SIZE 0.16 BY 0.16 ;
END MAS1561

MACRO MAS1562
   SIZE 0.16 BY 0.16 ;
END MAS1562

MACRO MAS1563
   SIZE 0.16 BY 0.16 ;
END MAS1563

MACRO MAS1564
   SIZE 0.16 BY 0.16 ;
END MAS1564

MACRO MAS1565
   SIZE 0.16 BY 0.16 ;
END MAS1565

MACRO MAS1566
   SIZE 0.16 BY 0.16 ;
END MAS1566

MACRO MAS1567
   SIZE 0.16 BY 0.16 ;
END MAS1567

MACRO MAS1568
   SIZE 0.16 BY 0.16 ;
END MAS1568

MACRO MAS1569
   SIZE 0.16 BY 0.16 ;
END MAS1569

MACRO MAS1570
   SIZE 0.16 BY 0.16 ;
END MAS1570

MACRO MAS1571
   SIZE 0.16 BY 0.16 ;
END MAS1571

MACRO MAS1572
   SIZE 0.16 BY 0.16 ;
END MAS1572

MACRO MAS1573
   SIZE 0.16 BY 0.16 ;
END MAS1573

MACRO MAS1574
   SIZE 0.16 BY 0.16 ;
END MAS1574

MACRO MAS1575
   SIZE 0.16 BY 0.16 ;
END MAS1575

MACRO MAS1576
   SIZE 0.16 BY 0.16 ;
END MAS1576

MACRO MAS1577
   SIZE 0.16 BY 0.16 ;
END MAS1577

MACRO MAS1578
   SIZE 0.16 BY 0.16 ;
END MAS1578

MACRO MAS1579
   SIZE 0.16 BY 0.16 ;
END MAS1579

MACRO MAS1580
   SIZE 0.16 BY 0.16 ;
END MAS1580

MACRO MAS1581
   SIZE 0.16 BY 0.16 ;
END MAS1581

MACRO MAS1582
   SIZE 0.16 BY 0.16 ;
END MAS1582

MACRO MAS1583
   SIZE 0.16 BY 0.16 ;
END MAS1583

MACRO MAS1584
   SIZE 0.16 BY 0.16 ;
END MAS1584

MACRO MAS1585
   SIZE 0.16 BY 0.16 ;
END MAS1585

MACRO MAS1586
   SIZE 0.16 BY 0.16 ;
END MAS1586

MACRO MAS1587
   SIZE 0.16 BY 0.16 ;
END MAS1587

MACRO MAS1588
   SIZE 0.16 BY 0.16 ;
END MAS1588

MACRO MAS1589
   SIZE 0.16 BY 0.16 ;
END MAS1589

MACRO MAS1590
   SIZE 0.16 BY 0.16 ;
END MAS1590

MACRO MAS1591
   SIZE 0.16 BY 0.16 ;
END MAS1591

MACRO MAS1592
   SIZE 0.16 BY 0.16 ;
END MAS1592

MACRO MAS1593
   SIZE 0.16 BY 0.16 ;
END MAS1593

MACRO MAS1594
   SIZE 0.16 BY 0.16 ;
END MAS1594

MACRO MAS1595
   SIZE 0.16 BY 0.16 ;
END MAS1595

MACRO MAS1596
   SIZE 0.16 BY 0.16 ;
END MAS1596

MACRO MAS1597
   SIZE 0.16 BY 0.16 ;
END MAS1597

MACRO MAS1598
   SIZE 0.16 BY 0.16 ;
END MAS1598

MACRO MAS1599
   SIZE 0.16 BY 0.16 ;
END MAS1599

MACRO MAS1600
   SIZE 0.16 BY 0.16 ;
END MAS1600

MACRO MAS1601
   SIZE 0.16 BY 0.16 ;
END MAS1601

MACRO MAS1602
   SIZE 0.16 BY 0.16 ;
END MAS1602

MACRO MAS1603
   SIZE 0.16 BY 0.16 ;
END MAS1603

MACRO MAS1604
   SIZE 0.16 BY 0.16 ;
END MAS1604

MACRO MAS1605
   SIZE 0.16 BY 0.16 ;
END MAS1605

MACRO MAS1606
   SIZE 0.16 BY 0.16 ;
END MAS1606

MACRO MAS1607
   SIZE 0.16 BY 0.16 ;
END MAS1607

MACRO MAS1608
   SIZE 0.16 BY 0.16 ;
END MAS1608

MACRO MAS1609
   SIZE 0.16 BY 0.16 ;
END MAS1609

MACRO MAS1610
   SIZE 0.16 BY 0.16 ;
END MAS1610

MACRO MAS1611
   SIZE 0.16 BY 0.16 ;
END MAS1611

MACRO MAS1612
   SIZE 0.16 BY 0.16 ;
END MAS1612

MACRO MAS1613
   SIZE 0.16 BY 0.16 ;
END MAS1613

MACRO MAS1614
   SIZE 0.16 BY 0.16 ;
END MAS1614

MACRO MAS1615
   SIZE 0.16 BY 0.16 ;
END MAS1615

MACRO MAS1616
   SIZE 0.16 BY 0.16 ;
END MAS1616

MACRO MAS1617
   SIZE 0.16 BY 0.16 ;
END MAS1617

MACRO MAS1618
   SIZE 0.16 BY 0.16 ;
END MAS1618

MACRO MAS1619
   SIZE 0.16 BY 0.16 ;
END MAS1619

MACRO MAS1620
   SIZE 0.16 BY 0.16 ;
END MAS1620

MACRO MAS1621
   SIZE 0.16 BY 0.16 ;
END MAS1621

MACRO MAS1622
   SIZE 0.16 BY 0.16 ;
END MAS1622

MACRO MAS1623
   SIZE 0.16 BY 0.16 ;
END MAS1623

MACRO MAS1624
   SIZE 0.16 BY 0.16 ;
END MAS1624

MACRO MAS1625
   SIZE 0.16 BY 0.16 ;
END MAS1625

MACRO MAS1626
   SIZE 0.16 BY 0.16 ;
END MAS1626

MACRO MAS1627
   SIZE 0.16 BY 0.16 ;
END MAS1627

MACRO MAS1628
   SIZE 0.18 BY 0.16 ;
END MAS1628

MACRO MAS1629
   SIZE 0.18 BY 0.16 ;
END MAS1629

MACRO MAS1630
   SIZE 0.18 BY 0.16 ;
END MAS1630

MACRO MAS1631
   SIZE 0.18 BY 0.16 ;
END MAS1631

MACRO MAS1632
   SIZE 0.18 BY 0.16 ;
END MAS1632

MACRO MAS1633
   SIZE 0.18 BY 0.16 ;
END MAS1633

MACRO MAS1634
   SIZE 0.18 BY 0.16 ;
END MAS1634

MACRO MAS1635
   SIZE 0.18 BY 0.16 ;
END MAS1635

MACRO MAS1636
   SIZE 0.18 BY 0.16 ;
END MAS1636

MACRO MAS1637
   SIZE 0.18 BY 0.16 ;
END MAS1637

MACRO MAS1638
   SIZE 0.18 BY 0.16 ;
END MAS1638

MACRO MAS1639
   SIZE 0.18 BY 0.16 ;
END MAS1639

MACRO MAS1640
   SIZE 0.18 BY 0.16 ;
END MAS1640

MACRO MAS1641
   SIZE 0.18 BY 0.16 ;
END MAS1641

MACRO MAS1642
   SIZE 0.18 BY 0.16 ;
END MAS1642

MACRO MAS1643
   SIZE 0.18 BY 0.16 ;
END MAS1643

MACRO MAS1644
   SIZE 0.18 BY 0.16 ;
END MAS1644

MACRO MAS1645
   SIZE 0.18 BY 0.16 ;
END MAS1645

MACRO MAS1646
   SIZE 0.18 BY 0.16 ;
END MAS1646

MACRO MAS1647
   SIZE 0.18 BY 0.16 ;
END MAS1647

MACRO MAS1648
   SIZE 0.18 BY 0.16 ;
END MAS1648

MACRO MAS1649
   SIZE 0.18 BY 0.16 ;
END MAS1649

MACRO MAS1650
   SIZE 0.18 BY 0.16 ;
END MAS1650

MACRO MAS1651
   SIZE 0.18 BY 0.16 ;
END MAS1651

MACRO MAS1652
   SIZE 0.18 BY 0.16 ;
END MAS1652

MACRO MAS1653
   SIZE 0.18 BY 0.16 ;
END MAS1653

MACRO MAS1654
   SIZE 0.18 BY 0.16 ;
END MAS1654

MACRO MAS1655
   SIZE 0.18 BY 0.16 ;
END MAS1655

MACRO MAS1656
   SIZE 0.18 BY 0.16 ;
END MAS1656

MACRO MAS1657
   SIZE 0.18 BY 0.16 ;
END MAS1657

MACRO MAS1658
   SIZE 0.18 BY 0.16 ;
END MAS1658

MACRO MAS1659
   SIZE 0.18 BY 0.16 ;
END MAS1659

MACRO MAS1660
   SIZE 0.18 BY 0.16 ;
END MAS1660

MACRO MAS1661
   SIZE 0.18 BY 0.16 ;
END MAS1661

MACRO MAS1662
   SIZE 0.18 BY 0.16 ;
END MAS1662

MACRO MAS1663
   SIZE 0.18 BY 0.16 ;
END MAS1663

MACRO MAS1664
   SIZE 0.18 BY 0.16 ;
END MAS1664

MACRO MAS1665
   SIZE 0.18 BY 0.16 ;
END MAS1665

MACRO MAS1666
   SIZE 0.18 BY 0.16 ;
END MAS1666

MACRO MAS1667
   SIZE 0.18 BY 0.16 ;
END MAS1667

MACRO MAS1668
   SIZE 0.18 BY 0.16 ;
END MAS1668

MACRO MAS1669
   SIZE 0.18 BY 0.16 ;
END MAS1669

MACRO MAS1670
   SIZE 0.18 BY 0.16 ;
END MAS1670

MACRO MAS1671
   SIZE 0.18 BY 0.16 ;
END MAS1671

MACRO MAS1672
   SIZE 0.18 BY 0.16 ;
END MAS1672

MACRO MAS1673
   SIZE 0.18 BY 0.16 ;
END MAS1673

MACRO MAS1674
   SIZE 0.18 BY 0.16 ;
END MAS1674

MACRO MAS1675
   SIZE 0.18 BY 0.16 ;
END MAS1675

MACRO MAS1676
   SIZE 0.18 BY 0.16 ;
END MAS1676

MACRO MAS1677
   SIZE 0.18 BY 0.16 ;
END MAS1677

MACRO MAS1678
   SIZE 0.18 BY 0.16 ;
END MAS1678

MACRO MAS1679
   SIZE 0.18 BY 0.16 ;
END MAS1679

MACRO MAS1680
   SIZE 0.18 BY 0.16 ;
END MAS1680

MACRO MAS1681
   SIZE 0.18 BY 0.16 ;
END MAS1681

MACRO MAS1682
   SIZE 0.18 BY 0.16 ;
END MAS1682

MACRO MAS1683
   SIZE 0.18 BY 0.16 ;
END MAS1683

MACRO MAS1684
   SIZE 0.18 BY 0.16 ;
END MAS1684

MACRO MAS1685
   SIZE 0.18 BY 0.16 ;
END MAS1685

MACRO MAS1686
   SIZE 0.18 BY 0.16 ;
END MAS1686

MACRO MAS1687
   SIZE 0.18 BY 0.16 ;
END MAS1687

MACRO MAS1688
   SIZE 0.18 BY 0.16 ;
END MAS1688

MACRO MAS1689
   SIZE 0.18 BY 0.16 ;
END MAS1689

MACRO MAS1690
   SIZE 0.18 BY 0.16 ;
END MAS1690

MACRO MAS1691
   SIZE 0.18 BY 0.16 ;
END MAS1691

MACRO MAS1692
   SIZE 0.18 BY 0.16 ;
END MAS1692

MACRO MAS1693
   SIZE 0.18 BY 0.16 ;
END MAS1693

MACRO MAS1694
   SIZE 0.18 BY 0.16 ;
END MAS1694

MACRO MAS1695
   SIZE 0.18 BY 0.16 ;
END MAS1695

MACRO MAS1696
   SIZE 0.18 BY 0.16 ;
END MAS1696

MACRO MAS1697
   SIZE 0.18 BY 0.16 ;
END MAS1697

MACRO MAS1698
   SIZE 0.18 BY 0.16 ;
END MAS1698

MACRO MAS1699
   SIZE 0.18 BY 0.16 ;
END MAS1699

MACRO MAS1700
   SIZE 0.18 BY 0.16 ;
END MAS1700

MACRO MAS1701
   SIZE 0.18 BY 0.16 ;
END MAS1701

MACRO MAS1702
   SIZE 0.18 BY 0.16 ;
END MAS1702

MACRO MAS1703
   SIZE 0.18 BY 0.16 ;
END MAS1703

MACRO MAS1704
   SIZE 0.18 BY 0.16 ;
END MAS1704

MACRO MAS1705
   SIZE 0.18 BY 0.16 ;
END MAS1705

MACRO MAS1706
   SIZE 0.18 BY 0.16 ;
END MAS1706

MACRO MAS1707
   SIZE 0.18 BY 0.16 ;
END MAS1707

MACRO MAS1708
   SIZE 0.18 BY 0.16 ;
END MAS1708

MACRO MAS1709
   SIZE 0.18 BY 0.16 ;
END MAS1709

MACRO MAS1710
   SIZE 0.18 BY 0.16 ;
END MAS1710

MACRO MAS1711
   SIZE 0.18 BY 0.16 ;
END MAS1711

MACRO MAS1712
   SIZE 0.18 BY 0.16 ;
END MAS1712

MACRO MAS1713
   SIZE 0.18 BY 0.16 ;
END MAS1713

MACRO MAS1714
   SIZE 0.18 BY 0.16 ;
END MAS1714

MACRO MAS1715
   SIZE 0.18 BY 0.16 ;
END MAS1715

MACRO MAS1716
   SIZE 0.18 BY 0.16 ;
END MAS1716

MACRO MAS1717
   SIZE 0.18 BY 0.16 ;
END MAS1717

MACRO MAS1718
   SIZE 0.18 BY 0.16 ;
END MAS1718

MACRO MAS1719
   SIZE 0.18 BY 0.16 ;
END MAS1719

MACRO MAS1720
   SIZE 0.18 BY 0.16 ;
END MAS1720

MACRO MAS1721
   SIZE 0.18 BY 0.16 ;
END MAS1721

MACRO MAS1722
   SIZE 0.18 BY 0.16 ;
END MAS1722

MACRO MAS1723
   SIZE 0.18 BY 0.16 ;
END MAS1723

MACRO MAS1724
   SIZE 0.18 BY 0.16 ;
END MAS1724

MACRO MAS1725
   SIZE 0.18 BY 0.16 ;
END MAS1725

MACRO MAS1726
   SIZE 0.18 BY 0.16 ;
END MAS1726

MACRO MAS1727
   SIZE 0.18 BY 0.16 ;
END MAS1727

MACRO MAS1728
   SIZE 0.18 BY 0.16 ;
END MAS1728

MACRO MAS1729
   SIZE 0.18 BY 0.16 ;
END MAS1729

MACRO MAS1730
   SIZE 0.18 BY 0.16 ;
END MAS1730

MACRO MAS1731
   SIZE 0.18 BY 0.16 ;
END MAS1731

MACRO MAS1732
   SIZE 0.18 BY 0.16 ;
END MAS1732

MACRO MAS1733
   SIZE 0.18 BY 0.16 ;
END MAS1733

MACRO MAS1734
   SIZE 0.18 BY 0.16 ;
END MAS1734

MACRO MAS1735
   SIZE 0.18 BY 0.16 ;
END MAS1735

MACRO MAS1736
   SIZE 0.18 BY 0.16 ;
END MAS1736

MACRO MAS1737
   SIZE 0.18 BY 0.16 ;
END MAS1737

MACRO MAS1738
   SIZE 0.18 BY 0.16 ;
END MAS1738

MACRO MAS1739
   SIZE 0.18 BY 0.16 ;
END MAS1739

MACRO MAS1740
   SIZE 0.18 BY 0.16 ;
END MAS1740

MACRO MAS1741
   SIZE 0.18 BY 0.16 ;
END MAS1741

MACRO MAS1742
   SIZE 0.18 BY 0.16 ;
END MAS1742

MACRO MAS1743
   SIZE 0.18 BY 0.16 ;
END MAS1743

MACRO MAS1744
   SIZE 0.18 BY 0.16 ;
END MAS1744

MACRO MAS1745
   SIZE 0.18 BY 0.16 ;
END MAS1745

MACRO MAS1746
   SIZE 0.18 BY 0.16 ;
END MAS1746

MACRO MAS1747
   SIZE 0.18 BY 0.16 ;
END MAS1747

MACRO MAS1748
   SIZE 0.18 BY 0.16 ;
END MAS1748

MACRO MAS1749
   SIZE 0.18 BY 0.16 ;
END MAS1749

MACRO MAS1750
   SIZE 0.18 BY 0.16 ;
END MAS1750

MACRO MAS1751
   SIZE 0.18 BY 0.16 ;
END MAS1751

MACRO MAS1752
   SIZE 0.18 BY 0.16 ;
END MAS1752

MACRO MAS1753
   SIZE 0.18 BY 0.16 ;
END MAS1753

MACRO MAS1754
   SIZE 0.18 BY 0.16 ;
END MAS1754

MACRO MAS1755
   SIZE 0.18 BY 0.16 ;
END MAS1755

MACRO MAS1756
   SIZE 0.18 BY 0.16 ;
END MAS1756

MACRO MAS1757
   SIZE 0.18 BY 0.16 ;
END MAS1757

MACRO MAS1758
   SIZE 0.2 BY 0.16 ;
END MAS1758

MACRO MAS1759
   SIZE 0.2 BY 0.16 ;
END MAS1759

MACRO MAS1760
   SIZE 0.2 BY 0.16 ;
END MAS1760

MACRO MAS1761
   SIZE 0.2 BY 0.16 ;
END MAS1761

MACRO MAS1762
   SIZE 0.2 BY 0.16 ;
END MAS1762

MACRO MAS1763
   SIZE 0.2 BY 0.16 ;
END MAS1763

MACRO MAS1764
   SIZE 0.2 BY 0.16 ;
END MAS1764

MACRO MAS1765
   SIZE 0.2 BY 0.16 ;
END MAS1765

MACRO MAS1766
   SIZE 0.2 BY 0.16 ;
END MAS1766

MACRO MAS1767
   SIZE 0.2 BY 0.16 ;
END MAS1767

MACRO MAS1768
   SIZE 0.2 BY 0.16 ;
END MAS1768

MACRO MAS1769
   SIZE 0.2 BY 0.16 ;
END MAS1769

MACRO MAS1770
   SIZE 0.2 BY 0.16 ;
END MAS1770

MACRO MAS1771
   SIZE 0.2 BY 0.16 ;
END MAS1771

MACRO MAS1772
   SIZE 0.2 BY 0.16 ;
END MAS1772

MACRO MAS1773
   SIZE 0.2 BY 0.16 ;
END MAS1773

MACRO MAS1774
   SIZE 0.2 BY 0.16 ;
END MAS1774

MACRO MAS1775
   SIZE 0.2 BY 0.16 ;
END MAS1775

MACRO MAS1776
   SIZE 0.2 BY 0.16 ;
END MAS1776

MACRO MAS1777
   SIZE 0.2 BY 0.16 ;
END MAS1777

MACRO MAS1778
   SIZE 0.2 BY 0.16 ;
END MAS1778

MACRO MAS1779
   SIZE 0.2 BY 0.16 ;
END MAS1779

MACRO MAS1780
   SIZE 0.2 BY 0.16 ;
END MAS1780

MACRO MAS1781
   SIZE 0.2 BY 0.16 ;
END MAS1781

MACRO MAS1782
   SIZE 0.2 BY 0.16 ;
END MAS1782

MACRO MAS1783
   SIZE 0.2 BY 0.16 ;
END MAS1783

MACRO MAS1784
   SIZE 0.2 BY 0.16 ;
END MAS1784

MACRO MAS1785
   SIZE 0.2 BY 0.16 ;
END MAS1785

MACRO MAS1786
   SIZE 0.2 BY 0.16 ;
END MAS1786

MACRO MAS1787
   SIZE 0.2 BY 0.16 ;
END MAS1787

MACRO MAS1788
   SIZE 0.2 BY 0.16 ;
END MAS1788

MACRO MAS1789
   SIZE 0.2 BY 0.16 ;
END MAS1789

MACRO MAS1790
   SIZE 0.2 BY 0.16 ;
END MAS1790

MACRO MAS1791
   SIZE 0.2 BY 0.16 ;
END MAS1791

MACRO MAS1792
   SIZE 0.2 BY 0.16 ;
END MAS1792

MACRO MAS1793
   SIZE 0.2 BY 0.16 ;
END MAS1793

MACRO MAS1794
   SIZE 0.2 BY 0.16 ;
END MAS1794

MACRO MAS1795
   SIZE 0.2 BY 0.16 ;
END MAS1795

MACRO MAS1796
   SIZE 0.2 BY 0.16 ;
END MAS1796

MACRO MAS1797
   SIZE 0.2 BY 0.16 ;
END MAS1797

MACRO MAS1798
   SIZE 0.2 BY 0.16 ;
END MAS1798

MACRO MAS1799
   SIZE 0.2 BY 0.16 ;
END MAS1799

MACRO MAS1800
   SIZE 0.2 BY 0.16 ;
END MAS1800

MACRO MAS1801
   SIZE 0.2 BY 0.16 ;
END MAS1801

MACRO MAS1802
   SIZE 0.2 BY 0.16 ;
END MAS1802

MACRO MAS1803
   SIZE 0.2 BY 0.16 ;
END MAS1803

MACRO MAS1804
   SIZE 0.2 BY 0.16 ;
END MAS1804

MACRO MAS1805
   SIZE 0.2 BY 0.16 ;
END MAS1805

MACRO MAS1806
   SIZE 0.2 BY 0.16 ;
END MAS1806

MACRO MAS1807
   SIZE 0.2 BY 0.16 ;
END MAS1807

MACRO MAS1808
   SIZE 0.2 BY 0.16 ;
END MAS1808

MACRO MAS1809
   SIZE 0.2 BY 0.16 ;
END MAS1809

MACRO MAS1810
   SIZE 0.2 BY 0.16 ;
END MAS1810

MACRO MAS1811
   SIZE 0.2 BY 0.16 ;
END MAS1811

MACRO MAS1812
   SIZE 0.2 BY 0.16 ;
END MAS1812

MACRO MAS1813
   SIZE 0.2 BY 0.16 ;
END MAS1813

MACRO MAS1814
   SIZE 0.2 BY 0.16 ;
END MAS1814

MACRO MAS1815
   SIZE 0.2 BY 0.16 ;
END MAS1815

MACRO MAS1816
   SIZE 0.2 BY 0.16 ;
END MAS1816

MACRO MAS1817
   SIZE 0.2 BY 0.16 ;
END MAS1817

MACRO MAS1818
   SIZE 0.2 BY 0.16 ;
END MAS1818

MACRO MAS1819
   SIZE 0.2 BY 0.16 ;
END MAS1819

MACRO MAS1820
   SIZE 0.2 BY 0.16 ;
END MAS1820

MACRO MAS1821
   SIZE 0.2 BY 0.16 ;
END MAS1821

MACRO MAS1822
   SIZE 0.2 BY 0.16 ;
END MAS1822

MACRO MAS1823
   SIZE 0.2 BY 0.16 ;
END MAS1823

MACRO MAS1824
   SIZE 0.2 BY 0.16 ;
END MAS1824

MACRO MAS1825
   SIZE 0.2 BY 0.16 ;
END MAS1825

MACRO MAS1826
   SIZE 0.2 BY 0.16 ;
END MAS1826

MACRO MAS1827
   SIZE 0.2 BY 0.16 ;
END MAS1827

MACRO MAS1828
   SIZE 0.2 BY 0.16 ;
END MAS1828

MACRO MAS1829
   SIZE 0.2 BY 0.16 ;
END MAS1829

MACRO MAS1830
   SIZE 0.2 BY 0.16 ;
END MAS1830

MACRO MAS1831
   SIZE 0.2 BY 0.16 ;
END MAS1831

MACRO MAS1832
   SIZE 0.2 BY 0.16 ;
END MAS1832

MACRO MAS1833
   SIZE 0.2 BY 0.16 ;
END MAS1833

MACRO MAS1834
   SIZE 0.2 BY 0.16 ;
END MAS1834

MACRO MAS1835
   SIZE 0.2 BY 0.16 ;
END MAS1835

MACRO MAS1836
   SIZE 0.2 BY 0.16 ;
END MAS1836

MACRO MAS1837
   SIZE 0.2 BY 0.16 ;
END MAS1837

MACRO MAS1838
   SIZE 0.2 BY 0.16 ;
END MAS1838

MACRO MAS1839
   SIZE 0.2 BY 0.16 ;
END MAS1839

MACRO MAS1840
   SIZE 0.2 BY 0.16 ;
END MAS1840

MACRO MAS1841
   SIZE 0.2 BY 0.16 ;
END MAS1841

MACRO MAS1842
   SIZE 0.2 BY 0.16 ;
END MAS1842

MACRO MAS1843
   SIZE 0.2 BY 0.16 ;
END MAS1843

MACRO MAS1844
   SIZE 0.2 BY 0.16 ;
END MAS1844

MACRO MAS1845
   SIZE 0.2 BY 0.16 ;
END MAS1845

MACRO MAS1846
   SIZE 0.2 BY 0.16 ;
END MAS1846

MACRO MAS1847
   SIZE 0.2 BY 0.16 ;
END MAS1847

MACRO MAS1848
   SIZE 0.2 BY 0.16 ;
END MAS1848

MACRO MAS1849
   SIZE 0.2 BY 0.16 ;
END MAS1849

MACRO MAS1850
   SIZE 0.2 BY 0.16 ;
END MAS1850

MACRO MAS1851
   SIZE 0.2 BY 0.16 ;
END MAS1851

MACRO MAS1852
   SIZE 0.2 BY 0.16 ;
END MAS1852

MACRO MAS1853
   SIZE 0.2 BY 0.16 ;
END MAS1853

MACRO MAS1854
   SIZE 0.2 BY 0.16 ;
END MAS1854

MACRO MAS1855
   SIZE 0.2 BY 0.16 ;
END MAS1855

MACRO MAS1856
   SIZE 0.2 BY 0.16 ;
END MAS1856

MACRO MAS1857
   SIZE 0.2 BY 0.16 ;
END MAS1857

MACRO MAS1858
   SIZE 0.2 BY 0.16 ;
END MAS1858

MACRO MAS1859
   SIZE 0.2 BY 0.16 ;
END MAS1859

MACRO MAS1860
   SIZE 0.2 BY 0.16 ;
END MAS1860

MACRO MAS1861
   SIZE 0.2 BY 0.16 ;
END MAS1861

MACRO MAS1862
   SIZE 0.2 BY 0.16 ;
END MAS1862

MACRO MAS1863
   SIZE 0.2 BY 0.16 ;
END MAS1863

MACRO MAS1864
   SIZE 0.2 BY 0.16 ;
END MAS1864

MACRO MAS1865
   SIZE 0.2 BY 0.16 ;
END MAS1865

MACRO MAS1866
   SIZE 0.2 BY 0.16 ;
END MAS1866

MACRO MAS1867
   SIZE 0.2 BY 0.16 ;
END MAS1867

MACRO MAS1868
   SIZE 0.2 BY 0.16 ;
END MAS1868

MACRO MAS1869
   SIZE 0.2 BY 0.16 ;
END MAS1869

MACRO MAS1870
   SIZE 0.2 BY 0.16 ;
END MAS1870

MACRO MAS1871
   SIZE 0.2 BY 0.16 ;
END MAS1871

MACRO MAS1872
   SIZE 0.2 BY 0.16 ;
END MAS1872

MACRO MAS1873
   SIZE 0.2 BY 0.16 ;
END MAS1873

MACRO MAS1874
   SIZE 0.2 BY 0.16 ;
END MAS1874

MACRO MAS1875
   SIZE 0.2 BY 0.16 ;
END MAS1875

MACRO MAS1876
   SIZE 0.2 BY 0.16 ;
END MAS1876

MACRO MAS1877
   SIZE 0.2 BY 0.16 ;
END MAS1877

MACRO MAS1878
   SIZE 0.2 BY 0.16 ;
END MAS1878

MACRO MAS1879
   SIZE 0.2 BY 0.16 ;
END MAS1879

MACRO MAS1880
   SIZE 0.2 BY 0.16 ;
END MAS1880

MACRO MAS1881
   SIZE 0.2 BY 0.16 ;
END MAS1881

MACRO MAS1882
   SIZE 0.22 BY 0.16 ;
END MAS1882

MACRO MAS1883
   SIZE 0.22 BY 0.16 ;
END MAS1883

MACRO MAS1884
   SIZE 0.22 BY 0.16 ;
END MAS1884

MACRO MAS1885
   SIZE 0.22 BY 0.16 ;
END MAS1885

MACRO MAS1886
   SIZE 0.22 BY 0.16 ;
END MAS1886

MACRO MAS1887
   SIZE 0.22 BY 0.16 ;
END MAS1887

MACRO MAS1888
   SIZE 0.22 BY 0.16 ;
END MAS1888

MACRO MAS1889
   SIZE 0.22 BY 0.16 ;
END MAS1889

MACRO MAS1890
   SIZE 0.22 BY 0.16 ;
END MAS1890

MACRO MAS1891
   SIZE 0.22 BY 0.16 ;
END MAS1891

MACRO MAS1892
   SIZE 0.22 BY 0.16 ;
END MAS1892

MACRO MAS1893
   SIZE 0.22 BY 0.16 ;
END MAS1893

MACRO MAS1894
   SIZE 0.22 BY 0.16 ;
END MAS1894

MACRO MAS1895
   SIZE 0.22 BY 0.16 ;
END MAS1895

MACRO MAS1896
   SIZE 0.22 BY 0.16 ;
END MAS1896

MACRO MAS1897
   SIZE 0.22 BY 0.16 ;
END MAS1897

MACRO MAS1898
   SIZE 0.22 BY 0.16 ;
END MAS1898

MACRO MAS1899
   SIZE 0.22 BY 0.16 ;
END MAS1899

MACRO MAS1900
   SIZE 0.22 BY 0.16 ;
END MAS1900

MACRO MAS1901
   SIZE 0.22 BY 0.16 ;
END MAS1901

MACRO MAS1902
   SIZE 0.22 BY 0.16 ;
END MAS1902

MACRO MAS1903
   SIZE 0.22 BY 0.16 ;
END MAS1903

MACRO MAS1904
   SIZE 0.24 BY 0.16 ;
END MAS1904

MACRO MAS1905
   SIZE 0.24 BY 0.16 ;
END MAS1905

MACRO MAS1906
   SIZE 0.24 BY 0.16 ;
END MAS1906

MACRO MAS1907
   SIZE 0.24 BY 0.16 ;
END MAS1907

MACRO MAS1908
   SIZE 0.24 BY 0.16 ;
END MAS1908

MACRO MAS1909
   SIZE 0.24 BY 0.16 ;
END MAS1909

MACRO MAS1910
   SIZE 0.24 BY 0.16 ;
END MAS1910

MACRO MAS1911
   SIZE 0.24 BY 0.16 ;
END MAS1911

MACRO MAS1912
   SIZE 0.24 BY 0.16 ;
END MAS1912

MACRO MAS1913
   SIZE 0.24 BY 0.16 ;
END MAS1913

MACRO MAS1914
   SIZE 0.24 BY 0.16 ;
END MAS1914

MACRO MAS1915
   SIZE 0.24 BY 0.16 ;
END MAS1915

MACRO MAS1916
   SIZE 0.24 BY 0.16 ;
END MAS1916

MACRO MAS1917
   SIZE 0.24 BY 0.16 ;
END MAS1917

MACRO MAS1918
   SIZE 0.24 BY 0.16 ;
END MAS1918

MACRO MAS1919
   SIZE 0.24 BY 0.16 ;
END MAS1919

MACRO MAS1920
   SIZE 0.24 BY 0.16 ;
END MAS1920

MACRO MAS1921
   SIZE 0.24 BY 0.16 ;
END MAS1921

MACRO MAS1922
   SIZE 0.24 BY 0.16 ;
END MAS1922

MACRO MAS1923
   SIZE 0.24 BY 0.16 ;
END MAS1923

MACRO MAS1924
   SIZE 0.24 BY 0.16 ;
END MAS1924

MACRO MAS1925
   SIZE 0.24 BY 0.16 ;
END MAS1925

MACRO MAS1926
   SIZE 0.24 BY 0.16 ;
END MAS1926

MACRO MAS1927
   SIZE 0.24 BY 0.16 ;
END MAS1927

MACRO MAS1928
   SIZE 0.24 BY 0.16 ;
END MAS1928

MACRO MAS1929
   SIZE 0.24 BY 0.16 ;
END MAS1929

MACRO MAS1930
   SIZE 0.24 BY 0.16 ;
END MAS1930

MACRO MAS1931
   SIZE 0.24 BY 0.16 ;
END MAS1931

MACRO MAS1932
   SIZE 0.24 BY 0.16 ;
END MAS1932

MACRO MAS1933
   SIZE 0.24 BY 0.16 ;
END MAS1933

MACRO MAS1934
   SIZE 0.24 BY 0.16 ;
END MAS1934

MACRO MAS1935
   SIZE 0.24 BY 0.16 ;
END MAS1935

MACRO MAS1936
   SIZE 0.24 BY 0.16 ;
END MAS1936

MACRO MAS1937
   SIZE 0.24 BY 0.16 ;
END MAS1937

MACRO MAS1938
   SIZE 0.24 BY 0.16 ;
END MAS1938

MACRO MAS1939
   SIZE 0.24 BY 0.16 ;
END MAS1939

MACRO MAS1940
   SIZE 0.24 BY 0.16 ;
END MAS1940

MACRO MAS1941
   SIZE 0.24 BY 0.16 ;
END MAS1941

MACRO MAS1942
   SIZE 0.24 BY 0.16 ;
END MAS1942

MACRO MAS1943
   SIZE 0.24 BY 0.16 ;
END MAS1943

MACRO MAS1944
   SIZE 0.24 BY 0.16 ;
END MAS1944

MACRO MAS1945
   SIZE 0.24 BY 0.16 ;
END MAS1945

MACRO MAS1946
   SIZE 0.24 BY 0.16 ;
END MAS1946

MACRO MAS1947
   SIZE 0.24 BY 0.16 ;
END MAS1947

MACRO MAS1948
   SIZE 0.24 BY 0.16 ;
END MAS1948

MACRO MAS1949
   SIZE 0.24 BY 0.16 ;
END MAS1949

MACRO MAS1950
   SIZE 0.24 BY 0.16 ;
END MAS1950

MACRO MAS1951
   SIZE 0.24 BY 0.16 ;
END MAS1951

MACRO MAS1952
   SIZE 0.24 BY 0.16 ;
END MAS1952

MACRO MAS1953
   SIZE 0.24 BY 0.16 ;
END MAS1953

MACRO MAS1954
   SIZE 0.24 BY 0.16 ;
END MAS1954

MACRO MAS1955
   SIZE 0.24 BY 0.16 ;
END MAS1955

MACRO MAS1956
   SIZE 0.24 BY 0.16 ;
END MAS1956

MACRO MAS1957
   SIZE 0.24 BY 0.16 ;
END MAS1957

MACRO MAS1958
   SIZE 0.24 BY 0.16 ;
END MAS1958

MACRO MAS1959
   SIZE 0.24 BY 0.16 ;
END MAS1959

MACRO MAS1960
   SIZE 0.24 BY 0.16 ;
END MAS1960

MACRO MAS1961
   SIZE 0.24 BY 0.16 ;
END MAS1961

MACRO MAS1962
   SIZE 0.24 BY 0.16 ;
END MAS1962

MACRO MAS1963
   SIZE 0.24 BY 0.16 ;
END MAS1963

MACRO MAS1964
   SIZE 0.24 BY 0.16 ;
END MAS1964

MACRO MAS1965
   SIZE 0.24 BY 0.16 ;
END MAS1965

MACRO MAS1966
   SIZE 0.24 BY 0.16 ;
END MAS1966

MACRO MAS1967
   SIZE 0.24 BY 0.16 ;
END MAS1967

MACRO MAS1968
   SIZE 0.24 BY 0.16 ;
END MAS1968

MACRO MAS1969
   SIZE 0.24 BY 0.16 ;
END MAS1969

MACRO MAS1970
   SIZE 0.24 BY 0.16 ;
END MAS1970

MACRO MAS1971
   SIZE 0.24 BY 0.16 ;
END MAS1971

MACRO MAS1972
   SIZE 0.24 BY 0.16 ;
END MAS1972

MACRO MAS1973
   SIZE 0.24 BY 0.16 ;
END MAS1973

MACRO MAS1974
   SIZE 0.24 BY 0.16 ;
END MAS1974

MACRO MAS1975
   SIZE 0.24 BY 0.16 ;
END MAS1975

MACRO MAS1976
   SIZE 0.24 BY 0.16 ;
END MAS1976

MACRO MAS1977
   SIZE 0.24 BY 0.16 ;
END MAS1977

MACRO MAS1978
   SIZE 0.24 BY 0.16 ;
END MAS1978

MACRO MAS1979
   SIZE 0.24 BY 0.16 ;
END MAS1979

MACRO MAS1980
   SIZE 0.24 BY 0.16 ;
END MAS1980

MACRO MAS1981
   SIZE 0.24 BY 0.16 ;
END MAS1981

MACRO MAS1982
   SIZE 0.24 BY 0.16 ;
END MAS1982

MACRO MAS1983
   SIZE 0.24 BY 0.16 ;
END MAS1983

MACRO MAS1984
   SIZE 0.24 BY 0.16 ;
END MAS1984

MACRO MAS1985
   SIZE 0.24 BY 0.16 ;
END MAS1985

MACRO MAS1986
   SIZE 0.24 BY 0.16 ;
END MAS1986

MACRO MAS1987
   SIZE 0.24 BY 0.16 ;
END MAS1987

MACRO MAS1988
   SIZE 0.24 BY 0.16 ;
END MAS1988

MACRO MAS1989
   SIZE 0.24 BY 0.16 ;
END MAS1989

MACRO MAS1990
   SIZE 0.24 BY 0.16 ;
END MAS1990

MACRO MAS1991
   SIZE 0.24 BY 0.16 ;
END MAS1991

MACRO MAS1992
   SIZE 0.24 BY 0.16 ;
END MAS1992

MACRO MAS1993
   SIZE 0.24 BY 0.16 ;
END MAS1993

MACRO MAS1994
   SIZE 0.24 BY 0.16 ;
END MAS1994

MACRO MAS1995
   SIZE 0.24 BY 0.16 ;
END MAS1995

MACRO MAS1996
   SIZE 0.24 BY 0.16 ;
END MAS1996

MACRO MAS1997
   SIZE 0.24 BY 0.16 ;
END MAS1997

MACRO MAS1998
   SIZE 0.24 BY 0.16 ;
END MAS1998

MACRO MAS1999
   SIZE 0.24 BY 0.16 ;
END MAS1999

MACRO MAS2000
   SIZE 0.24 BY 0.16 ;
END MAS2000

MACRO MAS2001
   SIZE 0.24 BY 0.16 ;
END MAS2001

MACRO MAS2002
   SIZE 0.24 BY 0.16 ;
END MAS2002

MACRO MAS2003
   SIZE 0.24 BY 0.16 ;
END MAS2003

MACRO MAS2004
   SIZE 0.24 BY 0.16 ;
END MAS2004

MACRO MAS2005
   SIZE 0.24 BY 0.16 ;
END MAS2005

MACRO MAS2006
   SIZE 0.24 BY 0.16 ;
END MAS2006

MACRO MAS2007
   SIZE 0.24 BY 0.16 ;
END MAS2007

MACRO MAS2008
   SIZE 0.24 BY 0.16 ;
END MAS2008

MACRO MAS2009
   SIZE 0.24 BY 0.16 ;
END MAS2009

MACRO MAS2010
   SIZE 0.24 BY 0.16 ;
END MAS2010

MACRO MAS2011
   SIZE 0.24 BY 0.16 ;
END MAS2011

MACRO MAS2012
   SIZE 0.24 BY 0.16 ;
END MAS2012

MACRO MAS2013
   SIZE 0.24 BY 0.16 ;
END MAS2013

MACRO MAS2014
   SIZE 0.24 BY 0.16 ;
END MAS2014

MACRO MAS2015
   SIZE 0.24 BY 0.16 ;
END MAS2015

MACRO MAS2016
   SIZE 0.24 BY 0.16 ;
END MAS2016

MACRO MAS2017
   SIZE 0.24 BY 0.16 ;
END MAS2017

MACRO MAS2018
   SIZE 0.24 BY 0.16 ;
END MAS2018

MACRO MAS2019
   SIZE 0.24 BY 0.16 ;
END MAS2019

MACRO MAS2020
   SIZE 0.24 BY 0.16 ;
END MAS2020

MACRO MAS2021
   SIZE 0.24 BY 0.16 ;
END MAS2021

MACRO MAS2022
   SIZE 0.24 BY 0.16 ;
END MAS2022

MACRO MAS2023
   SIZE 0.24 BY 0.16 ;
END MAS2023

MACRO MAS2024
   SIZE 0.24 BY 0.16 ;
END MAS2024

MACRO MAS2025
   SIZE 0.24 BY 0.16 ;
END MAS2025

MACRO MAS2026
   SIZE 0.24 BY 0.16 ;
END MAS2026

MACRO MAS2027
   SIZE 0.24 BY 0.16 ;
END MAS2027

MACRO MAS2028
   SIZE 0.24 BY 0.16 ;
END MAS2028

MACRO MAS2029
   SIZE 0.24 BY 0.16 ;
END MAS2029

MACRO MAS2030
   SIZE 0.24 BY 0.16 ;
END MAS2030

MACRO MAS2031
   SIZE 0.24 BY 0.16 ;
END MAS2031

MACRO MAS2032
   SIZE 0.24 BY 0.16 ;
END MAS2032

MACRO MAS2033
   SIZE 0.24 BY 0.16 ;
END MAS2033

MACRO MAS2034
   SIZE 0.24 BY 0.16 ;
END MAS2034

MACRO MAS2035
   SIZE 0.24 BY 0.16 ;
END MAS2035

MACRO MAS2036
   SIZE 0.24 BY 0.16 ;
END MAS2036

MACRO MAS2037
   SIZE 0.24 BY 0.16 ;
END MAS2037

MACRO MAS2038
   SIZE 0.24 BY 0.16 ;
END MAS2038

MACRO MAS2039
   SIZE 0.24 BY 0.16 ;
END MAS2039

MACRO MAS2040
   SIZE 0.24 BY 0.16 ;
END MAS2040

MACRO MAS2041
   SIZE 0.24 BY 0.16 ;
END MAS2041

MACRO MAS2042
   SIZE 0.24 BY 0.16 ;
END MAS2042

MACRO MAS2043
   SIZE 0.24 BY 0.16 ;
END MAS2043

MACRO MAS2044
   SIZE 0.24 BY 0.16 ;
END MAS2044

MACRO MAS2045
   SIZE 0.24 BY 0.16 ;
END MAS2045

MACRO MAS2046
   SIZE 0.24 BY 0.16 ;
END MAS2046

MACRO MAS2047
   SIZE 0.24 BY 0.16 ;
END MAS2047

MACRO MAS2048
   SIZE 0.24 BY 0.16 ;
END MAS2048

MACRO MAS2049
   SIZE 0.24 BY 0.16 ;
END MAS2049

MACRO MAS2050
   SIZE 0.24 BY 0.16 ;
END MAS2050

MACRO MAS2051
   SIZE 0.24 BY 0.16 ;
END MAS2051

MACRO MAS2052
   SIZE 0.24 BY 0.16 ;
END MAS2052

MACRO MAS2053
   SIZE 0.24 BY 0.16 ;
END MAS2053

MACRO MAS2054
   SIZE 0.24 BY 0.16 ;
END MAS2054

MACRO MAS2055
   SIZE 0.24 BY 0.16 ;
END MAS2055

MACRO MAS2056
   SIZE 0.24 BY 0.16 ;
END MAS2056

MACRO MAS2057
   SIZE 0.24 BY 0.16 ;
END MAS2057

MACRO MAS2058
   SIZE 0.24 BY 0.16 ;
END MAS2058

MACRO MAS2059
   SIZE 0.24 BY 0.16 ;
END MAS2059

MACRO MAS2060
   SIZE 0.24 BY 0.16 ;
END MAS2060

MACRO MAS2061
   SIZE 0.24 BY 0.16 ;
END MAS2061

MACRO MAS2062
   SIZE 0.24 BY 0.16 ;
END MAS2062

MACRO MAS2063
   SIZE 0.24 BY 0.16 ;
END MAS2063

MACRO MAS2064
   SIZE 0.24 BY 0.16 ;
END MAS2064

MACRO MAS2065
   SIZE 0.24 BY 0.16 ;
END MAS2065

MACRO MAS2066
   SIZE 0.24 BY 0.16 ;
END MAS2066

MACRO MAS2067
   SIZE 0.24 BY 0.16 ;
END MAS2067

MACRO MAS2068
   SIZE 0.24 BY 0.16 ;
END MAS2068

MACRO MAS2069
   SIZE 0.24 BY 0.16 ;
END MAS2069

MACRO MAS2070
   SIZE 0.24 BY 0.16 ;
END MAS2070

MACRO MAS2071
   SIZE 0.24 BY 0.16 ;
END MAS2071

MACRO MAS2072
   SIZE 0.24 BY 0.16 ;
END MAS2072

MACRO MAS2073
   SIZE 0.24 BY 0.16 ;
END MAS2073

MACRO MAS2074
   SIZE 0.24 BY 0.16 ;
END MAS2074

MACRO MAS2075
   SIZE 0.24 BY 0.16 ;
END MAS2075

MACRO MAS2076
   SIZE 0.24 BY 0.16 ;
END MAS2076

MACRO MAS2077
   SIZE 0.24 BY 0.16 ;
END MAS2077

MACRO MAS2078
   SIZE 0.24 BY 0.16 ;
END MAS2078

MACRO MAS2079
   SIZE 0.24 BY 0.16 ;
END MAS2079

MACRO MAS2080
   SIZE 0.24 BY 0.16 ;
END MAS2080

MACRO MAS2081
   SIZE 0.24 BY 0.16 ;
END MAS2081

MACRO MAS2082
   SIZE 0.24 BY 0.16 ;
END MAS2082

MACRO MAS2083
   SIZE 0.24 BY 0.16 ;
END MAS2083

MACRO MAS2084
   SIZE 0.24 BY 0.16 ;
END MAS2084

MACRO MAS2085
   SIZE 0.24 BY 0.16 ;
END MAS2085

MACRO MAS2086
   SIZE 0.24 BY 0.16 ;
END MAS2086

MACRO MAS2087
   SIZE 0.24 BY 0.16 ;
END MAS2087

MACRO MAS2088
   SIZE 0.24 BY 0.16 ;
END MAS2088

MACRO MAS2089
   SIZE 0.24 BY 0.16 ;
END MAS2089

MACRO MAS2090
   SIZE 0.24 BY 0.16 ;
END MAS2090

MACRO MAS2091
   SIZE 0.24 BY 0.16 ;
END MAS2091

MACRO MAS2092
   SIZE 0.24 BY 0.16 ;
END MAS2092

MACRO MAS2093
   SIZE 0.24 BY 0.16 ;
END MAS2093

MACRO MAS2094
   SIZE 0.24 BY 0.16 ;
END MAS2094

MACRO MAS2095
   SIZE 0.24 BY 0.16 ;
END MAS2095

MACRO MAS2096
   SIZE 0.24 BY 0.16 ;
END MAS2096

MACRO MAS2097
   SIZE 0.24 BY 0.16 ;
END MAS2097

MACRO MAS2098
   SIZE 0.24 BY 0.16 ;
END MAS2098

MACRO MAS2099
   SIZE 0.24 BY 0.16 ;
END MAS2099

MACRO MAS2100
   SIZE 0.24 BY 0.16 ;
END MAS2100

MACRO MAS2101
   SIZE 0.24 BY 0.16 ;
END MAS2101

MACRO MAS2102
   SIZE 0.24 BY 0.16 ;
END MAS2102

MACRO MAS2103
   SIZE 0.24 BY 0.16 ;
END MAS2103

MACRO MAS2104
   SIZE 0.24 BY 0.16 ;
END MAS2104

MACRO MAS2105
   SIZE 0.24 BY 0.16 ;
END MAS2105

MACRO MAS2106
   SIZE 0.24 BY 0.16 ;
END MAS2106

MACRO MAS2107
   SIZE 0.24 BY 0.16 ;
END MAS2107

MACRO MAS2108
   SIZE 0.24 BY 0.16 ;
END MAS2108

MACRO MAS2109
   SIZE 0.24 BY 0.16 ;
END MAS2109

MACRO MAS2110
   SIZE 0.24 BY 0.16 ;
END MAS2110

MACRO MAS2111
   SIZE 0.24 BY 0.16 ;
END MAS2111

MACRO MAS2112
   SIZE 0.24 BY 0.16 ;
END MAS2112

MACRO MAS2113
   SIZE 0.24 BY 0.16 ;
END MAS2113

MACRO MAS2114
   SIZE 0.24 BY 0.16 ;
END MAS2114

MACRO MAS2115
   SIZE 0.24 BY 0.16 ;
END MAS2115

MACRO MAS2116
   SIZE 0.24 BY 0.16 ;
END MAS2116

MACRO MAS2117
   SIZE 0.24 BY 0.16 ;
END MAS2117

MACRO MAS2118
   SIZE 0.24 BY 0.16 ;
END MAS2118

MACRO MAS2119
   SIZE 0.24 BY 0.16 ;
END MAS2119

MACRO MAS2120
   SIZE 0.24 BY 0.16 ;
END MAS2120

MACRO MAS2121
   SIZE 0.24 BY 0.16 ;
END MAS2121

MACRO MAS2122
   SIZE 0.24 BY 0.16 ;
END MAS2122

MACRO MAS2123
   SIZE 0.24 BY 0.16 ;
END MAS2123

MACRO MAS2124
   SIZE 0.24 BY 0.16 ;
END MAS2124

MACRO MAS2125
   SIZE 0.24 BY 0.16 ;
END MAS2125

MACRO MAS2126
   SIZE 0.24 BY 0.16 ;
END MAS2126

MACRO MAS2127
   SIZE 0.24 BY 0.16 ;
END MAS2127

MACRO MAS2128
   SIZE 0.24 BY 0.16 ;
END MAS2128

MACRO MAS2129
   SIZE 0.24 BY 0.16 ;
END MAS2129

MACRO MAS2130
   SIZE 0.24 BY 0.16 ;
END MAS2130

MACRO MAS2131
   SIZE 0.24 BY 0.16 ;
END MAS2131

MACRO MAS2132
   SIZE 0.24 BY 0.16 ;
END MAS2132

MACRO MAS2133
   SIZE 0.24 BY 0.16 ;
END MAS2133

MACRO MAS2134
   SIZE 0.24 BY 0.16 ;
END MAS2134

MACRO MAS2135
   SIZE 0.24 BY 0.16 ;
END MAS2135

MACRO MAS2136
   SIZE 0.24 BY 0.16 ;
END MAS2136

MACRO MAS2137
   SIZE 0.24 BY 0.16 ;
END MAS2137

MACRO MAS2138
   SIZE 0.24 BY 0.16 ;
END MAS2138

MACRO MAS2139
   SIZE 0.24 BY 0.16 ;
END MAS2139

MACRO MAS2140
   SIZE 0.24 BY 0.16 ;
END MAS2140

MACRO MAS2141
   SIZE 0.24 BY 0.16 ;
END MAS2141

MACRO MAS2142
   SIZE 0.24 BY 0.16 ;
END MAS2142

MACRO MAS2143
   SIZE 0.24 BY 0.16 ;
END MAS2143

MACRO MAS2144
   SIZE 0.24 BY 0.16 ;
END MAS2144

MACRO MAS2145
   SIZE 0.24 BY 0.16 ;
END MAS2145

MACRO MAS2146
   SIZE 0.24 BY 0.16 ;
END MAS2146

MACRO MAS2147
   SIZE 0.24 BY 0.16 ;
END MAS2147

MACRO MAS2148
   SIZE 0.24 BY 0.16 ;
END MAS2148

MACRO MAS2149
   SIZE 0.24 BY 0.16 ;
END MAS2149

MACRO MAS2150
   SIZE 0.24 BY 0.16 ;
END MAS2150

MACRO MAS2151
   SIZE 0.24 BY 0.16 ;
END MAS2151

MACRO MAS2152
   SIZE 0.24 BY 0.16 ;
END MAS2152

MACRO MAS2153
   SIZE 0.24 BY 0.16 ;
END MAS2153

MACRO MAS2154
   SIZE 0.26 BY 0.16 ;
END MAS2154

MACRO MAS2155
   SIZE 0.26 BY 0.16 ;
END MAS2155

MACRO MAS2156
   SIZE 0.26 BY 0.16 ;
END MAS2156

MACRO MAS2157
   SIZE 0.26 BY 0.16 ;
END MAS2157

MACRO MAS2158
   SIZE 0.26 BY 0.16 ;
END MAS2158

MACRO MAS2159
   SIZE 0.26 BY 0.16 ;
END MAS2159

MACRO MAS2160
   SIZE 0.26 BY 0.16 ;
END MAS2160

MACRO MAS2161
   SIZE 0.26 BY 0.16 ;
END MAS2161

MACRO MAS2162
   SIZE 0.26 BY 0.16 ;
END MAS2162

MACRO MAS2163
   SIZE 0.26 BY 0.16 ;
END MAS2163

MACRO MAS2164
   SIZE 0.26 BY 0.16 ;
END MAS2164

MACRO MAS2165
   SIZE 0.26 BY 0.16 ;
END MAS2165

MACRO MAS2166
   SIZE 0.26 BY 0.16 ;
END MAS2166

MACRO MAS2167
   SIZE 0.26 BY 0.16 ;
END MAS2167

MACRO MAS2168
   SIZE 0.26 BY 0.16 ;
END MAS2168

MACRO MAS2169
   SIZE 0.26 BY 0.16 ;
END MAS2169

MACRO MAS2170
   SIZE 0.26 BY 0.16 ;
END MAS2170

MACRO MAS2171
   SIZE 0.26 BY 0.16 ;
END MAS2171

MACRO MAS2172
   SIZE 0.26 BY 0.16 ;
END MAS2172

MACRO MAS2173
   SIZE 0.26 BY 0.16 ;
END MAS2173

MACRO MAS2174
   SIZE 0.26 BY 0.16 ;
END MAS2174

MACRO MAS2175
   SIZE 0.26 BY 0.16 ;
END MAS2175

MACRO MAS2176
   SIZE 0.26 BY 0.16 ;
END MAS2176

MACRO MAS2177
   SIZE 0.26 BY 0.16 ;
END MAS2177

MACRO MAS2178
   SIZE 0.26 BY 0.16 ;
END MAS2178

MACRO MAS2179
   SIZE 0.26 BY 0.16 ;
END MAS2179

MACRO MAS2180
   SIZE 0.26 BY 0.16 ;
END MAS2180

MACRO MAS2181
   SIZE 0.26 BY 0.16 ;
END MAS2181

MACRO MAS2182
   SIZE 0.26 BY 0.16 ;
END MAS2182

MACRO MAS2183
   SIZE 0.26 BY 0.16 ;
END MAS2183

MACRO MAS2184
   SIZE 0.26 BY 0.16 ;
END MAS2184

MACRO MAS2185
   SIZE 0.26 BY 0.16 ;
END MAS2185

MACRO MAS2186
   SIZE 0.26 BY 0.16 ;
END MAS2186

MACRO MAS2187
   SIZE 0.26 BY 0.16 ;
END MAS2187

MACRO MAS2188
   SIZE 0.26 BY 0.16 ;
END MAS2188

MACRO MAS2189
   SIZE 0.26 BY 0.16 ;
END MAS2189

MACRO MAS2190
   SIZE 0.26 BY 0.16 ;
END MAS2190

MACRO MAS2191
   SIZE 0.26 BY 0.16 ;
END MAS2191

MACRO MAS2192
   SIZE 0.26 BY 0.16 ;
END MAS2192

MACRO MAS2193
   SIZE 0.26 BY 0.16 ;
END MAS2193

MACRO MAS2194
   SIZE 0.26 BY 0.16 ;
END MAS2194

MACRO MAS2195
   SIZE 0.26 BY 0.16 ;
END MAS2195

MACRO MAS2196
   SIZE 0.26 BY 0.16 ;
END MAS2196

MACRO MAS2197
   SIZE 0.26 BY 0.16 ;
END MAS2197

MACRO MAS2198
   SIZE 0.26 BY 0.16 ;
END MAS2198

MACRO MAS2199
   SIZE 0.26 BY 0.16 ;
END MAS2199

MACRO MAS2200
   SIZE 0.26 BY 0.16 ;
END MAS2200

MACRO MAS2201
   SIZE 0.26 BY 0.16 ;
END MAS2201

MACRO MAS2202
   SIZE 0.26 BY 0.16 ;
END MAS2202

MACRO MAS2203
   SIZE 0.26 BY 0.16 ;
END MAS2203

MACRO MAS2204
   SIZE 0.26 BY 0.16 ;
END MAS2204

MACRO MAS2205
   SIZE 0.26 BY 0.16 ;
END MAS2205

MACRO MAS2206
   SIZE 0.26 BY 0.16 ;
END MAS2206

MACRO MAS2207
   SIZE 0.26 BY 0.16 ;
END MAS2207

MACRO MAS2208
   SIZE 0.26 BY 0.16 ;
END MAS2208

MACRO MAS2209
   SIZE 0.26 BY 0.16 ;
END MAS2209

MACRO MAS2210
   SIZE 0.26 BY 0.16 ;
END MAS2210

MACRO MAS2211
   SIZE 0.26 BY 0.16 ;
END MAS2211

MACRO MAS2212
   SIZE 0.26 BY 0.16 ;
END MAS2212

MACRO MAS2213
   SIZE 0.26 BY 0.16 ;
END MAS2213

MACRO MAS2214
   SIZE 0.26 BY 0.16 ;
END MAS2214

MACRO MAS2215
   SIZE 0.26 BY 0.16 ;
END MAS2215

MACRO MAS2216
   SIZE 0.26 BY 0.16 ;
END MAS2216

MACRO MAS2217
   SIZE 0.26 BY 0.16 ;
END MAS2217

MACRO MAS2218
   SIZE 0.26 BY 0.16 ;
END MAS2218

MACRO MAS2219
   SIZE 0.26 BY 0.16 ;
END MAS2219

MACRO MAS2220
   SIZE 0.26 BY 0.16 ;
END MAS2220

MACRO MAS2221
   SIZE 0.26 BY 0.16 ;
END MAS2221

MACRO MAS2222
   SIZE 0.26 BY 0.16 ;
END MAS2222

MACRO MAS2223
   SIZE 0.26 BY 0.16 ;
END MAS2223

MACRO MAS2224
   SIZE 0.26 BY 0.16 ;
END MAS2224

MACRO MAS2225
   SIZE 0.26 BY 0.16 ;
END MAS2225

MACRO MAS2226
   SIZE 0.26 BY 0.16 ;
END MAS2226

MACRO MAS2227
   SIZE 0.26 BY 0.16 ;
END MAS2227

MACRO MAS2228
   SIZE 0.28 BY 0.16 ;
END MAS2228

MACRO MAS2229
   SIZE 0.28 BY 0.16 ;
END MAS2229

MACRO MAS2230
   SIZE 0.28 BY 0.16 ;
END MAS2230

MACRO MAS2231
   SIZE 0.28 BY 0.16 ;
END MAS2231

MACRO MAS2232
   SIZE 0.28 BY 0.16 ;
END MAS2232

MACRO MAS2233
   SIZE 0.28 BY 0.16 ;
END MAS2233

MACRO MAS2234
   SIZE 0.28 BY 0.16 ;
END MAS2234

MACRO MAS2235
   SIZE 0.28 BY 0.16 ;
END MAS2235

MACRO MAS2236
   SIZE 0.28 BY 0.16 ;
END MAS2236

MACRO MAS2237
   SIZE 0.28 BY 0.16 ;
END MAS2237

MACRO MAS2238
   SIZE 0.28 BY 0.16 ;
END MAS2238

MACRO MAS2239
   SIZE 0.28 BY 0.16 ;
END MAS2239

MACRO MAS2240
   SIZE 0.28 BY 0.16 ;
END MAS2240

MACRO MAS2241
   SIZE 0.28 BY 0.16 ;
END MAS2241

MACRO MAS2242
   SIZE 0.28 BY 0.16 ;
END MAS2242

MACRO MAS2243
   SIZE 0.28 BY 0.16 ;
END MAS2243

MACRO MAS2244
   SIZE 0.28 BY 0.16 ;
END MAS2244

MACRO MAS2245
   SIZE 0.28 BY 0.16 ;
END MAS2245

MACRO MAS2246
   SIZE 0.28 BY 0.16 ;
END MAS2246

MACRO MAS2247
   SIZE 0.28 BY 0.16 ;
END MAS2247

MACRO MAS2248
   SIZE 0.28 BY 0.16 ;
END MAS2248

MACRO MAS2249
   SIZE 0.28 BY 0.16 ;
END MAS2249

MACRO MAS2250
   SIZE 0.28 BY 0.16 ;
END MAS2250

MACRO MAS2251
   SIZE 0.28 BY 0.16 ;
END MAS2251

MACRO MAS2252
   SIZE 0.28 BY 0.16 ;
END MAS2252

MACRO MAS2253
   SIZE 0.28 BY 0.16 ;
END MAS2253

MACRO MAS2254
   SIZE 0.28 BY 0.16 ;
END MAS2254

MACRO MAS2255
   SIZE 0.28 BY 0.16 ;
END MAS2255

MACRO MAS2256
   SIZE 0.28 BY 0.16 ;
END MAS2256

MACRO MAS2257
   SIZE 0.28 BY 0.16 ;
END MAS2257

MACRO MAS2258
   SIZE 0.28 BY 0.16 ;
END MAS2258

MACRO MAS2259
   SIZE 0.28 BY 0.16 ;
END MAS2259

MACRO MAS2260
   SIZE 0.28 BY 0.16 ;
END MAS2260

MACRO MAS2261
   SIZE 0.28 BY 0.16 ;
END MAS2261

MACRO MAS2262
   SIZE 0.28 BY 0.16 ;
END MAS2262

MACRO MAS2263
   SIZE 0.28 BY 0.16 ;
END MAS2263

MACRO MAS2264
   SIZE 0.28 BY 0.16 ;
END MAS2264

MACRO MAS2265
   SIZE 0.28 BY 0.16 ;
END MAS2265

MACRO MAS2266
   SIZE 0.28 BY 0.16 ;
END MAS2266

MACRO MAS2267
   SIZE 0.28 BY 0.16 ;
END MAS2267

MACRO MAS2268
   SIZE 0.28 BY 0.16 ;
END MAS2268

MACRO MAS2269
   SIZE 0.28 BY 0.16 ;
END MAS2269

MACRO MAS2270
   SIZE 0.28 BY 0.16 ;
END MAS2270

MACRO MAS2271
   SIZE 0.28 BY 0.16 ;
END MAS2271

MACRO MAS2272
   SIZE 0.28 BY 0.16 ;
END MAS2272

MACRO MAS2273
   SIZE 0.28 BY 0.16 ;
END MAS2273

MACRO MAS2274
   SIZE 0.28 BY 0.16 ;
END MAS2274

MACRO MAS2275
   SIZE 0.28 BY 0.16 ;
END MAS2275

MACRO MAS2276
   SIZE 0.28 BY 0.16 ;
END MAS2276

MACRO MAS2277
   SIZE 0.28 BY 0.16 ;
END MAS2277

MACRO MAS2278
   SIZE 0.28 BY 0.16 ;
END MAS2278

MACRO MAS2279
   SIZE 0.28 BY 0.16 ;
END MAS2279

MACRO MAS2280
   SIZE 0.28 BY 0.16 ;
END MAS2280

MACRO MAS2281
   SIZE 0.28 BY 0.16 ;
END MAS2281

MACRO MAS2282
   SIZE 0.28 BY 0.16 ;
END MAS2282

MACRO MAS2283
   SIZE 0.28 BY 0.16 ;
END MAS2283

MACRO MAS2284
   SIZE 0.28 BY 0.16 ;
END MAS2284

MACRO MAS2285
   SIZE 0.28 BY 0.16 ;
END MAS2285

MACRO MAS2286
   SIZE 0.28 BY 0.16 ;
END MAS2286

MACRO MAS2287
   SIZE 0.28 BY 0.16 ;
END MAS2287

MACRO MAS2288
   SIZE 0.28 BY 0.16 ;
END MAS2288

MACRO MAS2289
   SIZE 0.28 BY 0.16 ;
END MAS2289

MACRO MAS2290
   SIZE 0.28 BY 0.16 ;
END MAS2290

MACRO MAS2291
   SIZE 0.28 BY 0.16 ;
END MAS2291

MACRO MAS2292
   SIZE 0.28 BY 0.16 ;
END MAS2292

MACRO MAS2293
   SIZE 0.28 BY 0.16 ;
END MAS2293

MACRO MAS2294
   SIZE 0.28 BY 0.16 ;
END MAS2294

MACRO MAS2295
   SIZE 0.28 BY 0.16 ;
END MAS2295

MACRO MAS2296
   SIZE 0.28 BY 0.16 ;
END MAS2296

MACRO MAS2297
   SIZE 0.28 BY 0.16 ;
END MAS2297

MACRO MAS2298
   SIZE 0.28 BY 0.16 ;
END MAS2298

MACRO MAS2299
   SIZE 0.28 BY 0.16 ;
END MAS2299

MACRO MAS2300
   SIZE 0.28 BY 0.16 ;
END MAS2300

MACRO MAS2301
   SIZE 0.28 BY 0.16 ;
END MAS2301

MACRO MAS2302
   SIZE 0.28 BY 0.16 ;
END MAS2302

MACRO MAS2303
   SIZE 0.28 BY 0.16 ;
END MAS2303

MACRO MAS2304
   SIZE 0.28 BY 0.16 ;
END MAS2304

MACRO MAS2305
   SIZE 0.28 BY 0.16 ;
END MAS2305

MACRO MAS2306
   SIZE 0.28 BY 0.16 ;
END MAS2306

MACRO MAS2307
   SIZE 0.28 BY 0.16 ;
END MAS2307

MACRO MAS2308
   SIZE 0.28 BY 0.16 ;
END MAS2308

MACRO MAS2309
   SIZE 0.28 BY 0.16 ;
END MAS2309

MACRO MAS2310
   SIZE 0.28 BY 0.16 ;
END MAS2310

MACRO MAS2311
   SIZE 0.28 BY 0.16 ;
END MAS2311

MACRO MAS2312
   SIZE 0.28 BY 0.16 ;
END MAS2312

MACRO MAS2313
   SIZE 0.28 BY 0.16 ;
END MAS2313

MACRO MAS2314
   SIZE 0.28 BY 0.16 ;
END MAS2314

MACRO MAS2315
   SIZE 0.28 BY 0.16 ;
END MAS2315

MACRO MAS2316
   SIZE 0.28 BY 0.16 ;
END MAS2316

MACRO MAS2317
   SIZE 0.28 BY 0.16 ;
END MAS2317

MACRO MAS2318
   SIZE 0.28 BY 0.16 ;
END MAS2318

MACRO MAS2319
   SIZE 0.28 BY 0.16 ;
END MAS2319

MACRO MAS2320
   SIZE 0.28 BY 0.16 ;
END MAS2320

MACRO MAS2321
   SIZE 0.28 BY 0.16 ;
END MAS2321

MACRO MAS2322
   SIZE 0.28 BY 0.16 ;
END MAS2322

MACRO MAS2323
   SIZE 0.28 BY 0.16 ;
END MAS2323

MACRO MAS2324
   SIZE 0.28 BY 0.16 ;
END MAS2324

MACRO MAS2325
   SIZE 0.28 BY 0.16 ;
END MAS2325

MACRO MAS2326
   SIZE 0.28 BY 0.16 ;
END MAS2326

MACRO MAS2327
   SIZE 0.28 BY 0.16 ;
END MAS2327

MACRO MAS2328
   SIZE 0.28 BY 0.16 ;
END MAS2328

MACRO MAS2329
   SIZE 0.28 BY 0.16 ;
END MAS2329

MACRO MAS2330
   SIZE 0.28 BY 0.16 ;
END MAS2330

MACRO MAS2331
   SIZE 0.28 BY 0.16 ;
END MAS2331

MACRO MAS2332
   SIZE 0.28 BY 0.16 ;
END MAS2332

MACRO MAS2333
   SIZE 0.28 BY 0.16 ;
END MAS2333

MACRO MAS2334
   SIZE 0.28 BY 0.16 ;
END MAS2334

MACRO MAS2335
   SIZE 0.28 BY 0.16 ;
END MAS2335

MACRO MAS2336
   SIZE 0.28 BY 0.16 ;
END MAS2336

MACRO MAS2337
   SIZE 0.28 BY 0.16 ;
END MAS2337

MACRO MAS2338
   SIZE 0.28 BY 0.16 ;
END MAS2338

MACRO MAS2339
   SIZE 0.28 BY 0.16 ;
END MAS2339

MACRO MAS2340
   SIZE 0.28 BY 0.16 ;
END MAS2340

MACRO MAS2341
   SIZE 0.28 BY 0.16 ;
END MAS2341

MACRO MAS2342
   SIZE 0.3 BY 0.16 ;
END MAS2342

MACRO MAS2343
   SIZE 0.3 BY 0.16 ;
END MAS2343

MACRO MAS2344
   SIZE 0.3 BY 0.16 ;
END MAS2344

MACRO MAS2345
   SIZE 0.3 BY 0.16 ;
END MAS2345

MACRO MAS2346
   SIZE 0.3 BY 0.16 ;
END MAS2346

MACRO MAS2347
   SIZE 0.3 BY 0.16 ;
END MAS2347

MACRO MAS2348
   SIZE 0.3 BY 0.16 ;
END MAS2348

MACRO MAS2349
   SIZE 0.3 BY 0.16 ;
END MAS2349

MACRO MAS2350
   SIZE 0.3 BY 0.16 ;
END MAS2350

MACRO MAS2351
   SIZE 0.3 BY 0.16 ;
END MAS2351

MACRO MAS2352
   SIZE 0.3 BY 0.16 ;
END MAS2352

MACRO MAS2353
   SIZE 0.3 BY 0.16 ;
END MAS2353

MACRO MAS2354
   SIZE 0.3 BY 0.16 ;
END MAS2354

MACRO MAS2355
   SIZE 0.3 BY 0.16 ;
END MAS2355

MACRO MAS2356
   SIZE 0.3 BY 0.16 ;
END MAS2356

MACRO MAS2357
   SIZE 0.3 BY 0.16 ;
END MAS2357

MACRO MAS2358
   SIZE 0.3 BY 0.16 ;
END MAS2358

MACRO MAS2359
   SIZE 0.3 BY 0.16 ;
END MAS2359

MACRO MAS2360
   SIZE 0.3 BY 0.16 ;
END MAS2360

MACRO MAS2361
   SIZE 0.3 BY 0.16 ;
END MAS2361

MACRO MAS2362
   SIZE 0.3 BY 0.16 ;
END MAS2362

MACRO MAS2363
   SIZE 0.3 BY 0.16 ;
END MAS2363

MACRO MAS2364
   SIZE 0.3 BY 0.16 ;
END MAS2364

MACRO MAS2365
   SIZE 0.3 BY 0.16 ;
END MAS2365

MACRO MAS2366
   SIZE 0.3 BY 0.16 ;
END MAS2366

MACRO MAS2367
   SIZE 0.3 BY 0.16 ;
END MAS2367

MACRO MAS2368
   SIZE 0.3 BY 0.16 ;
END MAS2368

MACRO MAS2369
   SIZE 0.3 BY 0.16 ;
END MAS2369

MACRO MAS2370
   SIZE 0.3 BY 0.16 ;
END MAS2370

MACRO MAS2371
   SIZE 0.34 BY 0.16 ;
END MAS2371

MACRO MAS2372
   SIZE 0.34 BY 0.16 ;
END MAS2372

MACRO MAS2373
   SIZE 0.34 BY 0.16 ;
END MAS2373

MACRO MAS2374
   SIZE 0.34 BY 0.16 ;
END MAS2374

MACRO MAS2375
   SIZE 0.34 BY 0.16 ;
END MAS2375

MACRO MAS2376
   SIZE 0.34 BY 0.16 ;
END MAS2376

MACRO MAS2377
   SIZE 0.42 BY 0.16 ;
END MAS2377

MACRO MAS2378
   SIZE 0.42 BY 0.16 ;
END MAS2378

MACRO MAS2379
   SIZE 0.42 BY 0.16 ;
END MAS2379

MACRO MAS2380
   SIZE 0.42 BY 0.16 ;
END MAS2380

MACRO MAS2381
   SIZE 0.42 BY 0.16 ;
END MAS2381

MACRO MAS2382
   SIZE 0.42 BY 0.16 ;
END MAS2382

MACRO MAS2383
   SIZE 0.42 BY 0.16 ;
END MAS2383

MACRO MAS2384
   SIZE 0.42 BY 0.16 ;
END MAS2384

MACRO MAS2385
   SIZE 0.42 BY 0.16 ;
END MAS2385

MACRO MAS2386
   SIZE 0.42 BY 0.16 ;
END MAS2386

MACRO MAS2387
   SIZE 0.42 BY 0.16 ;
END MAS2387

MACRO MAS2388
   SIZE 0.42 BY 0.16 ;
END MAS2388

MACRO MAS2389
   SIZE 0.42 BY 0.16 ;
END MAS2389

MACRO MAS2390
   SIZE 0.42 BY 0.16 ;
END MAS2390

MACRO MAS2391
   SIZE 0.42 BY 0.16 ;
END MAS2391

MACRO MAS2392
   SIZE 0.42 BY 0.16 ;
END MAS2392

MACRO MAS2393
   SIZE 0.42 BY 0.16 ;
END MAS2393

MACRO MAS2394
   SIZE 0.42 BY 0.16 ;
END MAS2394

MACRO MAS2395
   SIZE 0.42 BY 0.16 ;
END MAS2395

MACRO MAS2396
   SIZE 0.42 BY 0.16 ;
END MAS2396

MACRO MAS2397
   SIZE 0.42 BY 0.16 ;
END MAS2397

MACRO MAS2398
   SIZE 0.42 BY 0.16 ;
END MAS2398

MACRO MAS2399
   SIZE 0.42 BY 0.16 ;
END MAS2399

MACRO MAS2400
   SIZE 0.42 BY 0.16 ;
END MAS2400

MACRO MAS2401
   SIZE 0.42 BY 0.16 ;
END MAS2401

MACRO MAS2402
   SIZE 0.42 BY 0.16 ;
END MAS2402

MACRO MAS2403
   SIZE 0.42 BY 0.16 ;
END MAS2403

MACRO MAS2404
   SIZE 0.42 BY 0.16 ;
END MAS2404

MACRO MAS2405
   SIZE 0.42 BY 0.16 ;
END MAS2405

MACRO MAS2406
   SIZE 0.42 BY 0.16 ;
END MAS2406

MACRO MAS2407
   SIZE 0.42 BY 0.16 ;
END MAS2407

MACRO MAS2408
   SIZE 0.42 BY 0.16 ;
END MAS2408

MACRO MAS2409
   SIZE 0.42 BY 0.16 ;
END MAS2409

MACRO MAS2410
   SIZE 0.42 BY 0.16 ;
END MAS2410

MACRO MAS2411
   SIZE 0.42 BY 0.16 ;
END MAS2411

MACRO MAS2412
   SIZE 0.42 BY 0.16 ;
END MAS2412

MACRO MAS2413
   SIZE 0.42 BY 0.16 ;
END MAS2413

MACRO MAS2414
   SIZE 0.42 BY 0.16 ;
END MAS2414

MACRO MAS2415
   SIZE 0.42 BY 0.16 ;
END MAS2415

MACRO MAS2416
   SIZE 0.42 BY 0.16 ;
END MAS2416

MACRO MAS2417
   SIZE 0.42 BY 0.16 ;
END MAS2417

MACRO MAS2418
   SIZE 0.42 BY 0.16 ;
END MAS2418

MACRO MAS2419
   SIZE 0.42 BY 0.16 ;
END MAS2419

MACRO MAS2420
   SIZE 0.42 BY 0.16 ;
END MAS2420

MACRO MAS2421
   SIZE 0.42 BY 0.16 ;
END MAS2421

MACRO MAS2422
   SIZE 0.42 BY 0.16 ;
END MAS2422

MACRO MAS2423
   SIZE 0.42 BY 0.16 ;
END MAS2423

MACRO MAS2424
   SIZE 0.42 BY 0.16 ;
END MAS2424

MACRO MAS2425
   SIZE 0.42 BY 0.16 ;
END MAS2425

MACRO MAS2426
   SIZE 0.42 BY 0.16 ;
END MAS2426

MACRO MAS2427
   SIZE 0.42 BY 0.16 ;
END MAS2427

MACRO MAS2428
   SIZE 0.42 BY 0.16 ;
END MAS2428

MACRO MAS2429
   SIZE 0.42 BY 0.16 ;
END MAS2429

MACRO MAS2430
   SIZE 0.42 BY 0.16 ;
END MAS2430

MACRO MAS2431
   SIZE 0.42 BY 0.16 ;
END MAS2431

MACRO MAS2432
   SIZE 0.42 BY 0.16 ;
END MAS2432

MACRO MAS2433
   SIZE 0.42 BY 0.16 ;
END MAS2433

MACRO MAS2434
   SIZE 0.42 BY 0.16 ;
END MAS2434

MACRO MAS2435
   SIZE 0.42 BY 0.16 ;
END MAS2435

MACRO MAS2436
   SIZE 0.42 BY 0.16 ;
END MAS2436

MACRO MAS2437
   SIZE 0.42 BY 0.16 ;
END MAS2437

MACRO MAS2438
   SIZE 0.42 BY 0.16 ;
END MAS2438

MACRO MAS2439
   SIZE 0.42 BY 0.16 ;
END MAS2439

MACRO MAS2440
   SIZE 0.42 BY 0.16 ;
END MAS2440

MACRO MAS2441
   SIZE 0.42 BY 0.16 ;
END MAS2441

MACRO MAS2442
   SIZE 0.42 BY 0.16 ;
END MAS2442

MACRO MAS2443
   SIZE 0.42 BY 0.16 ;
END MAS2443

MACRO MAS2444
   SIZE 0.42 BY 0.16 ;
END MAS2444

MACRO MAS2445
   SIZE 0.42 BY 0.16 ;
END MAS2445

MACRO MAS2446
   SIZE 0.42 BY 0.16 ;
END MAS2446

MACRO MAS2447
   SIZE 0.42 BY 0.16 ;
END MAS2447

MACRO MAS2448
   SIZE 0.42 BY 0.16 ;
END MAS2448

MACRO MAS2449
   SIZE 0.42 BY 0.16 ;
END MAS2449

MACRO MAS2450
   SIZE 0.42 BY 0.16 ;
END MAS2450

MACRO MAS2451
   SIZE 0.42 BY 0.16 ;
END MAS2451

MACRO MAS2452
   SIZE 0.42 BY 0.16 ;
END MAS2452

MACRO MAS2453
   SIZE 0.42 BY 0.16 ;
END MAS2453

MACRO MAS2454
   SIZE 0.42 BY 0.16 ;
END MAS2454

MACRO MAS2455
   SIZE 0.42 BY 0.16 ;
END MAS2455

MACRO MAS2456
   SIZE 0.42 BY 0.16 ;
END MAS2456

MACRO MAS2457
   SIZE 0.42 BY 0.16 ;
END MAS2457

MACRO MAS2458
   SIZE 0.42 BY 0.16 ;
END MAS2458

MACRO MAS2459
   SIZE 0.42 BY 0.16 ;
END MAS2459

MACRO MAS2460
   SIZE 0.42 BY 0.16 ;
END MAS2460

MACRO MAS2461
   SIZE 0.42 BY 0.16 ;
END MAS2461

MACRO MAS2462
   SIZE 0.42 BY 0.16 ;
END MAS2462

MACRO MAS2463
   SIZE 0.42 BY 0.16 ;
END MAS2463

MACRO MAS2464
   SIZE 0.42 BY 0.16 ;
END MAS2464

MACRO MAS2465
   SIZE 0.42 BY 0.16 ;
END MAS2465

MACRO MAS2466
   SIZE 0.42 BY 0.16 ;
END MAS2466

MACRO MAS2467
   SIZE 0.42 BY 0.16 ;
END MAS2467

MACRO MAS2468
   SIZE 0.42 BY 0.16 ;
END MAS2468

MACRO MAS2469
   SIZE 0.42 BY 0.16 ;
END MAS2469

MACRO MAS2470
   SIZE 0.42 BY 0.16 ;
END MAS2470

MACRO MAS2471
   SIZE 0.42 BY 0.16 ;
END MAS2471

MACRO MAS2472
   SIZE 0.42 BY 0.16 ;
END MAS2472

MACRO MAS2473
   SIZE 0.42 BY 0.16 ;
END MAS2473

MACRO MAS2474
   SIZE 0.42 BY 0.16 ;
END MAS2474

MACRO MAS2475
   SIZE 0.42 BY 0.16 ;
END MAS2475

MACRO MAS2476
   SIZE 0.42 BY 0.16 ;
END MAS2476

MACRO MAS2477
   SIZE 0.42 BY 0.16 ;
END MAS2477

MACRO MAS2478
   SIZE 0.42 BY 0.16 ;
END MAS2478

MACRO MAS2479
   SIZE 0.42 BY 0.16 ;
END MAS2479

MACRO MAS2480
   SIZE 0.42 BY 0.16 ;
END MAS2480

MACRO MAS2481
   SIZE 0.42 BY 0.16 ;
END MAS2481

MACRO MAS2482
   SIZE 0.42 BY 0.16 ;
END MAS2482

MACRO MAS2483
   SIZE 0.42 BY 0.16 ;
END MAS2483

MACRO MAS2484
   SIZE 0.42 BY 0.16 ;
END MAS2484

MACRO MAS2485
   SIZE 0.42 BY 0.16 ;
END MAS2485

MACRO MAS2486
   SIZE 0.42 BY 0.16 ;
END MAS2486

MACRO MAS2487
   SIZE 0.42 BY 0.16 ;
END MAS2487

MACRO MAS2488
   SIZE 0.42 BY 0.16 ;
END MAS2488

MACRO MAS2489
   SIZE 0.42 BY 0.16 ;
END MAS2489

MACRO MAS2490
   SIZE 0.42 BY 0.16 ;
END MAS2490

MACRO MAS2491
   SIZE 0.42 BY 0.16 ;
END MAS2491

MACRO MAS2492
   SIZE 0.42 BY 0.16 ;
END MAS2492

MACRO MAS2493
   SIZE 0.42 BY 0.16 ;
END MAS2493

MACRO MAS2494
   SIZE 0.42 BY 0.16 ;
END MAS2494

MACRO MAS2495
   SIZE 0.42 BY 0.16 ;
END MAS2495

MACRO MAS2496
   SIZE 0.42 BY 0.16 ;
END MAS2496

MACRO MAS2497
   SIZE 0.42 BY 0.16 ;
END MAS2497

MACRO MAS2498
   SIZE 0.42 BY 0.16 ;
END MAS2498

MACRO MAS2499
   SIZE 0.42 BY 0.16 ;
END MAS2499

MACRO MAS2500
   SIZE 0.42 BY 0.16 ;
END MAS2500

MACRO MAS2501
   SIZE 0.42 BY 0.16 ;
END MAS2501

MACRO MAS2502
   SIZE 0.42 BY 0.16 ;
END MAS2502

MACRO MAS2503
   SIZE 0.42 BY 0.16 ;
END MAS2503

MACRO MAS2504
   SIZE 0.42 BY 0.16 ;
END MAS2504

MACRO MAS2505
   SIZE 0.42 BY 0.16 ;
END MAS2505

MACRO MAS2506
   SIZE 0.42 BY 0.16 ;
END MAS2506

MACRO MAS2507
   SIZE 0.42 BY 0.16 ;
END MAS2507

MACRO MAS2508
   SIZE 0.42 BY 0.16 ;
END MAS2508

MACRO MAS2509
   SIZE 0.42 BY 0.16 ;
END MAS2509

MACRO MAS2510
   SIZE 0.42 BY 0.16 ;
END MAS2510

MACRO MAS2511
   SIZE 0.42 BY 0.16 ;
END MAS2511

MACRO MAS2512
   SIZE 0.42 BY 0.16 ;
END MAS2512

MACRO MAS2513
   SIZE 0.42 BY 0.16 ;
END MAS2513

MACRO MAS2514
   SIZE 0.42 BY 0.16 ;
END MAS2514

MACRO MAS2515
   SIZE 0.42 BY 0.16 ;
END MAS2515

MACRO MAS2516
   SIZE 0.42 BY 0.16 ;
END MAS2516

MACRO MAS2517
   SIZE 0.42 BY 0.16 ;
END MAS2517

MACRO MAS2518
   SIZE 0.42 BY 0.16 ;
END MAS2518

MACRO MAS2519
   SIZE 0.42 BY 0.16 ;
END MAS2519

MACRO MAS2520
   SIZE 0.42 BY 0.16 ;
END MAS2520

MACRO MAS2521
   SIZE 0.42 BY 0.16 ;
END MAS2521

MACRO MAS2522
   SIZE 0.42 BY 0.16 ;
END MAS2522

MACRO MAS2523
   SIZE 0.42 BY 0.16 ;
END MAS2523

MACRO MAS2524
   SIZE 0.42 BY 0.16 ;
END MAS2524

MACRO MAS2525
   SIZE 0.42 BY 0.16 ;
END MAS2525

MACRO MAS2526
   SIZE 0.42 BY 0.16 ;
END MAS2526

MACRO MAS2527
   SIZE 0.42 BY 0.16 ;
END MAS2527

MACRO MAS2528
   SIZE 0.42 BY 0.16 ;
END MAS2528

MACRO MAS2529
   SIZE 0.42 BY 0.16 ;
END MAS2529

MACRO MAS2530
   SIZE 0.42 BY 0.16 ;
END MAS2530

MACRO MAS2531
   SIZE 0.42 BY 0.16 ;
END MAS2531

MACRO MAS2532
   SIZE 0.42 BY 0.16 ;
END MAS2532

MACRO MAS2533
   SIZE 0.42 BY 0.16 ;
END MAS2533

MACRO MAS2534
   SIZE 0.42 BY 0.16 ;
END MAS2534

MACRO MAS2535
   SIZE 0.42 BY 0.16 ;
END MAS2535

MACRO MAS2536
   SIZE 0.42 BY 0.16 ;
END MAS2536

MACRO MAS2537
   SIZE 0.42 BY 0.16 ;
END MAS2537

MACRO MAS2538
   SIZE 0.42 BY 0.16 ;
END MAS2538

MACRO MAS2539
   SIZE 0.42 BY 0.16 ;
END MAS2539

MACRO MAS2540
   SIZE 0.42 BY 0.16 ;
END MAS2540

MACRO MAS2541
   SIZE 0.42 BY 0.16 ;
END MAS2541

MACRO MAS2542
   SIZE 0.42 BY 0.16 ;
END MAS2542

MACRO MAS2543
   SIZE 0.42 BY 0.16 ;
END MAS2543

MACRO MAS2544
   SIZE 0.42 BY 0.16 ;
END MAS2544

MACRO MAS2545
   SIZE 0.42 BY 0.16 ;
END MAS2545

MACRO MAS2546
   SIZE 0.42 BY 0.16 ;
END MAS2546

MACRO MAS2547
   SIZE 0.42 BY 0.16 ;
END MAS2547

MACRO MAS2548
   SIZE 0.42 BY 0.16 ;
END MAS2548

MACRO MAS2549
   SIZE 0.42 BY 0.16 ;
END MAS2549

MACRO MAS2550
   SIZE 0.42 BY 0.16 ;
END MAS2550

MACRO MAS2551
   SIZE 0.42 BY 0.16 ;
END MAS2551

MACRO MAS2552
   SIZE 0.42 BY 0.16 ;
END MAS2552

MACRO MAS2553
   SIZE 0.42 BY 0.16 ;
END MAS2553

MACRO MAS2554
   SIZE 0.42 BY 0.16 ;
END MAS2554

MACRO MAS2555
   SIZE 0.42 BY 0.16 ;
END MAS2555

MACRO MAS2556
   SIZE 0.42 BY 0.16 ;
END MAS2556

MACRO MAS2557
   SIZE 0.42 BY 0.16 ;
END MAS2557

MACRO MAS2558
   SIZE 0.42 BY 0.16 ;
END MAS2558

MACRO MAS2559
   SIZE 0.42 BY 0.16 ;
END MAS2559

MACRO MAS2560
   SIZE 0.42 BY 0.16 ;
END MAS2560

MACRO MAS2561
   SIZE 0.42 BY 0.16 ;
END MAS2561

MACRO MAS2562
   SIZE 0.42 BY 0.16 ;
END MAS2562

MACRO MAS2563
   SIZE 0.42 BY 0.16 ;
END MAS2563

MACRO MAS2564
   SIZE 0.42 BY 0.16 ;
END MAS2564

MACRO MAS2565
   SIZE 0.42 BY 0.16 ;
END MAS2565

MACRO MAS2566
   SIZE 0.42 BY 0.16 ;
END MAS2566

MACRO MAS2567
   SIZE 0.42 BY 0.16 ;
END MAS2567

MACRO MAS2568
   SIZE 0.42 BY 0.16 ;
END MAS2568

MACRO MAS2569
   SIZE 0.42 BY 0.16 ;
END MAS2569

MACRO MAS2570
   SIZE 0.42 BY 0.16 ;
END MAS2570

MACRO MAS2571
   SIZE 0.42 BY 0.16 ;
END MAS2571

MACRO MAS2572
   SIZE 0.42 BY 0.16 ;
END MAS2572

MACRO MAS2573
   SIZE 0.42 BY 0.16 ;
END MAS2573

MACRO MAS2574
   SIZE 0.42 BY 0.16 ;
END MAS2574

MACRO MAS2575
   SIZE 0.42 BY 0.16 ;
END MAS2575

MACRO MAS2576
   SIZE 0.42 BY 0.16 ;
END MAS2576

MACRO MAS2577
   SIZE 0.42 BY 0.16 ;
END MAS2577

MACRO MAS2578
   SIZE 0.42 BY 0.16 ;
END MAS2578

MACRO MAS2579
   SIZE 0.42 BY 0.16 ;
END MAS2579

MACRO MAS2580
   SIZE 0.42 BY 0.16 ;
END MAS2580

MACRO MAS2581
   SIZE 0.42 BY 0.16 ;
END MAS2581

MACRO MAS2582
   SIZE 0.42 BY 0.16 ;
END MAS2582

MACRO MAS2583
   SIZE 0.42 BY 0.16 ;
END MAS2583

MACRO MAS2584
   SIZE 0.42 BY 0.16 ;
END MAS2584

MACRO MAS2585
   SIZE 0.42 BY 0.16 ;
END MAS2585

MACRO MAS2586
   SIZE 0.42 BY 0.16 ;
END MAS2586

MACRO MAS2587
   SIZE 0.42 BY 0.16 ;
END MAS2587

MACRO MAS2588
   SIZE 0.42 BY 0.16 ;
END MAS2588

MACRO MAS2589
   SIZE 0.42 BY 0.16 ;
END MAS2589

MACRO MAS2590
   SIZE 0.42 BY 0.16 ;
END MAS2590

MACRO MAS2591
   SIZE 0.42 BY 0.16 ;
END MAS2591

MACRO MAS2592
   SIZE 0.42 BY 0.16 ;
END MAS2592

MACRO MAS2593
   SIZE 0.42 BY 0.16 ;
END MAS2593

MACRO MAS2594
   SIZE 0.42 BY 0.16 ;
END MAS2594

MACRO MAS2595
   SIZE 0.42 BY 0.16 ;
END MAS2595

MACRO MAS2596
   SIZE 0.42 BY 0.16 ;
END MAS2596

MACRO MAS2597
   SIZE 0.46 BY 0.16 ;
END MAS2597

MACRO MAS2598
   SIZE 0.46 BY 0.16 ;
END MAS2598

MACRO MAS2599
   SIZE 0.46 BY 0.16 ;
END MAS2599

MACRO MAS2600
   SIZE 0.63 BY 1.28 ;
END MAS2600

MACRO MAS2601
   SIZE 0.63 BY 1.28 ;
END MAS2601

MACRO MAS2602
   SIZE 0.63 BY 1.28 ;
END MAS2602

MACRO MAS2603
   SIZE 0.63 BY 1.28 ;
END MAS2603

MACRO MAS2604
   SIZE 0.63 BY 1.28 ;
END MAS2604

MACRO MAS2605
   SIZE 0.63 BY 1.28 ;
END MAS2605

MACRO MAS2606
   SIZE 0.63 BY 1.28 ;
END MAS2606

MACRO MAS2607
   SIZE 0.63 BY 1.28 ;
END MAS2607

MACRO MAS2608
   SIZE 0.63 BY 1.28 ;
END MAS2608

MACRO MAS2609
   SIZE 0.63 BY 1.28 ;
END MAS2609

MACRO MAS2610
   SIZE 0.63 BY 1.28 ;
END MAS2610

MACRO MAS2611
   SIZE 0.63 BY 1.28 ;
END MAS2611

MACRO MAS2612
   SIZE 0.63 BY 1.28 ;
END MAS2612

MACRO MAS2613
   SIZE 0.63 BY 1.28 ;
END MAS2613

MACRO MAS2614
   SIZE 0.63 BY 1.28 ;
END MAS2614

MACRO MAS2615
   SIZE 0.63 BY 1.28 ;
END MAS2615

MACRO MAS2616
   SIZE 0.63 BY 1.28 ;
END MAS2616

MACRO MAS2617
   SIZE 0.63 BY 1.28 ;
END MAS2617

MACRO MAS2618
   SIZE 0.63 BY 1.28 ;
END MAS2618

MACRO MAS2619
   SIZE 0.63 BY 1.28 ;
END MAS2619

MACRO MAS2620
   SIZE 0.63 BY 1.28 ;
END MAS2620

MACRO MAS2621
   SIZE 0.63 BY 1.28 ;
END MAS2621

MACRO MAS2622
   SIZE 0.63 BY 1.28 ;
END MAS2622

MACRO MAS2623
   SIZE 0.72 BY 1.12 ;
END MAS2623

MACRO MAS2624
   SIZE 0.72 BY 1.12 ;
END MAS2624

MACRO MAS2625
   SIZE 0.72 BY 1.12 ;
END MAS2625

MACRO MAS2626
   SIZE 0.72 BY 1.12 ;
END MAS2626

MACRO MAS2627
   SIZE 0.72 BY 1.12 ;
END MAS2627

MACRO MAS2628
   SIZE 0.72 BY 1.12 ;
END MAS2628

MACRO MAS2629
   SIZE 0.72 BY 1.12 ;
END MAS2629

MACRO MAS2630
   SIZE 0.72 BY 1.12 ;
END MAS2630

MACRO MAS2631
   SIZE 0.72 BY 1.12 ;
END MAS2631

MACRO MAS2632
   SIZE 0.72 BY 1.12 ;
END MAS2632

MACRO MAS2633
   SIZE 0.72 BY 1.12 ;
END MAS2633

MACRO MAS2634
   SIZE 0.72 BY 1.12 ;
END MAS2634

MACRO MAS2635
   SIZE 0.72 BY 1.12 ;
END MAS2635

MACRO MAS2636
   SIZE 0.72 BY 1.12 ;
END MAS2636

MACRO MAS2637
   SIZE 0.72 BY 1.12 ;
END MAS2637

MACRO MAS2638
   SIZE 0.72 BY 1.12 ;
END MAS2638

MACRO MAS2639
   SIZE 0.72 BY 1.12 ;
END MAS2639

MACRO MAS2640
   SIZE 0.72 BY 1.12 ;
END MAS2640

MACRO MAS2641
   SIZE 0.72 BY 1.12 ;
END MAS2641

MACRO MAS2642
   SIZE 0.72 BY 1.12 ;
END MAS2642

MACRO MAS2643
   SIZE 0.72 BY 1.12 ;
END MAS2643

MACRO MAS2644
   SIZE 0.72 BY 1.12 ;
END MAS2644

MACRO MAS2645
   SIZE 0.72 BY 1.12 ;
END MAS2645

MACRO MAS2646
   SIZE 0.72 BY 1.12 ;
END MAS2646

MACRO MAS2647
   SIZE 0.72 BY 1.12 ;
END MAS2647

MACRO MAS2648
   SIZE 0.72 BY 1.12 ;
END MAS2648

MACRO MAS2649
   SIZE 0.72 BY 1.12 ;
END MAS2649

MACRO MAS2650
   SIZE 0.72 BY 1.12 ;
END MAS2650

MACRO MAS2651
   SIZE 0.72 BY 1.12 ;
END MAS2651

MACRO MAS2652
   SIZE 0.72 BY 1.12 ;
END MAS2652

MACRO MAS2653
   SIZE 0.72 BY 1.12 ;
END MAS2653

MACRO MAS2654
   SIZE 0.72 BY 1.12 ;
END MAS2654

MACRO MAS2655
   SIZE 0.72 BY 1.12 ;
END MAS2655

MACRO MAS2656
   SIZE 0.72 BY 1.12 ;
END MAS2656

MACRO MAS2657
   SIZE 0.72 BY 1.12 ;
END MAS2657

MACRO MAS2658
   SIZE 0.84 BY 0.96 ;
END MAS2658

MACRO MAS2659
   SIZE 0.84 BY 0.96 ;
END MAS2659

MACRO MAS2660
   SIZE 0.84 BY 0.96 ;
END MAS2660

MACRO MAS2661
   SIZE 0.84 BY 0.96 ;
END MAS2661

MACRO MAS2662
   SIZE 0.84 BY 0.96 ;
END MAS2662

MACRO MAS2663
   SIZE 0.84 BY 0.96 ;
END MAS2663

MACRO MAS2664
   SIZE 0.84 BY 0.96 ;
END MAS2664

MACRO MAS2665
   SIZE 0.84 BY 0.96 ;
END MAS2665

MACRO MAS2666
   SIZE 0.84 BY 0.96 ;
END MAS2666

MACRO MAS2667
   SIZE 0.84 BY 0.96 ;
END MAS2667

MACRO MAS2668
   SIZE 0.84 BY 0.96 ;
END MAS2668

MACRO MAS2669
   SIZE 0.84 BY 0.96 ;
END MAS2669

MACRO MAS2670
   SIZE 0.84 BY 0.96 ;
END MAS2670

MACRO MAS2671
   SIZE 0.84 BY 0.96 ;
END MAS2671

MACRO MAS2672
   SIZE 0.84 BY 0.96 ;
END MAS2672

MACRO MAS2673
   SIZE 0.84 BY 0.96 ;
END MAS2673

MACRO MAS2674
   SIZE 0.84 BY 0.96 ;
END MAS2674

MACRO MAS2675
   SIZE 0.84 BY 0.96 ;
END MAS2675

MACRO MAS2676
   SIZE 0.84 BY 0.96 ;
END MAS2676

MACRO MAS2677
   SIZE 0.84 BY 0.96 ;
END MAS2677

MACRO MAS2678
   SIZE 0.84 BY 0.96 ;
END MAS2678

MACRO MAS2679
   SIZE 0.84 BY 0.96 ;
END MAS2679

MACRO MAS2680
   SIZE 0.84 BY 0.96 ;
END MAS2680

MACRO MAS2681
   SIZE 0.84 BY 0.96 ;
END MAS2681

MACRO MAS2682
   SIZE 0.84 BY 0.96 ;
END MAS2682

MACRO MAS2683
   SIZE 0.84 BY 0.96 ;
END MAS2683

MACRO MAS2684
   SIZE 0.84 BY 0.96 ;
END MAS2684

MACRO MAS2685
   SIZE 0.84 BY 0.96 ;
END MAS2685

MACRO MAS2686
   SIZE 0.84 BY 0.96 ;
END MAS2686

MACRO MAS2687
   SIZE 0.84 BY 0.96 ;
END MAS2687

MACRO MAS2688
   SIZE 0.84 BY 0.96 ;
END MAS2688

MACRO MAS2689
   SIZE 0.84 BY 0.96 ;
END MAS2689

MACRO MAS2690
   SIZE 0.84 BY 0.96 ;
END MAS2690

MACRO MAS2691
   SIZE 0.84 BY 0.96 ;
END MAS2691

MACRO MAS2692
   SIZE 0.84 BY 0.96 ;
END MAS2692

MACRO MAS2693
   SIZE 0.84 BY 0.96 ;
END MAS2693

MACRO MAS2694
   SIZE 0.84 BY 0.96 ;
END MAS2694

MACRO MAS2695
   SIZE 0.84 BY 0.96 ;
END MAS2695

MACRO MAS2696
   SIZE 0.84 BY 0.96 ;
END MAS2696

MACRO MAS2697
   SIZE 0.84 BY 0.96 ;
END MAS2697

MACRO MAS2698
   SIZE 0.84 BY 0.96 ;
END MAS2698

MACRO MAS2699
   SIZE 0.84 BY 0.96 ;
END MAS2699

MACRO MAS2700
   SIZE 0.84 BY 0.96 ;
END MAS2700

MACRO MAS2701
   SIZE 0.84 BY 0.96 ;
END MAS2701

MACRO MAS2702
   SIZE 0.84 BY 0.96 ;
END MAS2702

MACRO MAS2703
   SIZE 0.84 BY 0.96 ;
END MAS2703

MACRO MAS2704
   SIZE 0.84 BY 0.96 ;
END MAS2704

MACRO MAS2705
   SIZE 0.84 BY 0.96 ;
END MAS2705

MACRO MAS2706
   SIZE 0.84 BY 0.96 ;
END MAS2706

MACRO MAS2707
   SIZE 0.84 BY 0.96 ;
END MAS2707

MACRO MAS2708
   SIZE 0.84 BY 0.96 ;
END MAS2708

MACRO MAS2709
   SIZE 0.84 BY 0.96 ;
END MAS2709

MACRO MAS2710
   SIZE 0.84 BY 0.96 ;
END MAS2710

MACRO MAS2711
   SIZE 0.84 BY 0.96 ;
END MAS2711

MACRO MAS2712
   SIZE 0.84 BY 0.96 ;
END MAS2712

MACRO MAS2713
   SIZE 0.84 BY 0.96 ;
END MAS2713

MACRO MAS2714
   SIZE 0.84 BY 0.96 ;
END MAS2714

MACRO MAS2715
   SIZE 0.84 BY 0.96 ;
END MAS2715

MACRO MAS2716
   SIZE 0.84 BY 0.96 ;
END MAS2716

MACRO MAS2717
   SIZE 0.84 BY 0.96 ;
END MAS2717

MACRO MAS2718
   SIZE 0.84 BY 0.96 ;
END MAS2718

MACRO MAS2719
   SIZE 0.84 BY 0.96 ;
END MAS2719

MACRO MAS2720
   SIZE 0.84 BY 0.96 ;
END MAS2720

MACRO MAS2721
   SIZE 0.84 BY 0.96 ;
END MAS2721

MACRO MAS2722
   SIZE 0.84 BY 0.96 ;
END MAS2722

MACRO MAS2723
   SIZE 0.84 BY 0.96 ;
END MAS2723

MACRO MAS2724
   SIZE 1.26 BY 0.64 ;
END MAS2724

MACRO MAS2725
   SIZE 1.26 BY 0.64 ;
END MAS2725

MACRO MAS2726
   SIZE 1.01 BY 0.8 ;
END MAS2726

MACRO MAS2727
   SIZE 1.01 BY 0.8 ;
END MAS2727

MACRO MAS2728
   SIZE 1.01 BY 0.8 ;
END MAS2728

MACRO MAS2729
   SIZE 1.01 BY 0.8 ;
END MAS2729

MACRO MAS2730
   SIZE 1.01 BY 0.8 ;
END MAS2730

MACRO MAS2731
   SIZE 1.01 BY 0.8 ;
END MAS2731

MACRO MAS2732
   SIZE 1.01 BY 0.8 ;
END MAS2732

MACRO MAS2733
   SIZE 1.01 BY 0.8 ;
END MAS2733

MACRO MAS2734
   SIZE 1.01 BY 0.8 ;
END MAS2734

MACRO MAS2735
   SIZE 1.01 BY 0.8 ;
END MAS2735

MACRO MAS2736
   SIZE 1.01 BY 0.8 ;
END MAS2736

MACRO MAS2737
   SIZE 1.01 BY 0.8 ;
END MAS2737

MACRO MAS2738
   SIZE 1.01 BY 0.8 ;
END MAS2738

MACRO MAS2739
   SIZE 1.01 BY 0.8 ;
END MAS2739

MACRO MAS2740
   SIZE 1.01 BY 0.8 ;
END MAS2740

MACRO MAS2741
   SIZE 1.01 BY 0.8 ;
END MAS2741

MACRO MAS2742
   SIZE 1.01 BY 0.8 ;
END MAS2742

MACRO MAS2743
   SIZE 1.01 BY 0.8 ;
END MAS2743

MACRO MAS2744
   SIZE 1.01 BY 0.8 ;
END MAS2744

MACRO MAS2745
   SIZE 1.01 BY 0.8 ;
END MAS2745

MACRO MAS2746
   SIZE 1.01 BY 0.8 ;
END MAS2746

MACRO MAS2747
   SIZE 1.01 BY 0.8 ;
END MAS2747

MACRO MAS2748
   SIZE 1.01 BY 0.8 ;
END MAS2748

MACRO MAS2749
   SIZE 1.01 BY 0.8 ;
END MAS2749

MACRO MAS2750
   SIZE 1.01 BY 0.8 ;
END MAS2750

MACRO MAS2751
   SIZE 1.01 BY 0.8 ;
END MAS2751

MACRO MAS2752
   SIZE 1.01 BY 0.8 ;
END MAS2752

MACRO MAS2753
   SIZE 1.01 BY 0.8 ;
END MAS2753

MACRO MAS2754
   SIZE 1.01 BY 0.8 ;
END MAS2754

MACRO MAS2755
   SIZE 1.01 BY 0.8 ;
END MAS2755

MACRO MAS2756
   SIZE 1.01 BY 0.8 ;
END MAS2756

MACRO MAS2757
   SIZE 1.01 BY 0.8 ;
END MAS2757

MACRO MAS2758
   SIZE 1.01 BY 0.8 ;
END MAS2758

MACRO MAS2759
   SIZE 1.01 BY 0.8 ;
END MAS2759

MACRO MAS2760
   SIZE 1.01 BY 0.8 ;
END MAS2760

MACRO MAS2761
   SIZE 1.01 BY 0.8 ;
END MAS2761

MACRO MAS2762
   SIZE 1.01 BY 0.8 ;
END MAS2762

MACRO MAS2763
   SIZE 1.01 BY 0.8 ;
END MAS2763

MACRO MAS2764
   SIZE 1.01 BY 0.8 ;
END MAS2764

MACRO MAS2765
   SIZE 1.01 BY 0.8 ;
END MAS2765

MACRO MAS2766
   SIZE 1.01 BY 0.8 ;
END MAS2766

MACRO MAS2767
   SIZE 1.01 BY 0.8 ;
END MAS2767

MACRO MAS2768
   SIZE 1.01 BY 0.8 ;
END MAS2768

MACRO MAS2769
   SIZE 1.01 BY 0.8 ;
END MAS2769

MACRO MAS2770
   SIZE 1.01 BY 0.8 ;
END MAS2770

MACRO MAS2771
   SIZE 1.01 BY 0.8 ;
END MAS2771

MACRO MAS2772
   SIZE 1.01 BY 0.8 ;
END MAS2772

MACRO MAS2773
   SIZE 1.01 BY 0.8 ;
END MAS2773

MACRO MAS2774
   SIZE 1.01 BY 0.8 ;
END MAS2774

MACRO MAS2775
   SIZE 1.01 BY 0.8 ;
END MAS2775

MACRO MAS2776
   SIZE 1.01 BY 0.8 ;
END MAS2776

MACRO MAS2777
   SIZE 1.01 BY 0.8 ;
END MAS2777

MACRO MAS2778
   SIZE 1.01 BY 0.8 ;
END MAS2778

MACRO MAS2779
   SIZE 1.01 BY 0.8 ;
END MAS2779

MACRO MAS2780
   SIZE 1.01 BY 0.8 ;
END MAS2780

MACRO MAS2781
   SIZE 1.01 BY 0.8 ;
END MAS2781

MACRO MAS2782
   SIZE 1.01 BY 0.8 ;
END MAS2782

MACRO MAS2783
   SIZE 1.01 BY 0.8 ;
END MAS2783

MACRO MAS2784
   SIZE 1.01 BY 0.8 ;
END MAS2784

MACRO MAS2785
   SIZE 1.01 BY 0.8 ;
END MAS2785

MACRO MAS2786
   SIZE 1.01 BY 0.8 ;
END MAS2786

MACRO MAS2787
   SIZE 1.01 BY 0.8 ;
END MAS2787

MACRO MAS2788
   SIZE 1.01 BY 0.8 ;
END MAS2788

MACRO MAS2789
   SIZE 1.01 BY 0.8 ;
END MAS2789

MACRO MAS2790
   SIZE 1.01 BY 0.8 ;
END MAS2790

MACRO MAS2791
   SIZE 1.01 BY 0.8 ;
END MAS2791

MACRO MAS2792
   SIZE 1.01 BY 0.8 ;
END MAS2792

MACRO MAS2793
   SIZE 1.01 BY 0.8 ;
END MAS2793

MACRO MAS2794
   SIZE 1.01 BY 0.8 ;
END MAS2794

MACRO MAS2795
   SIZE 1.01 BY 0.8 ;
END MAS2795

MACRO MAS2796
   SIZE 1.01 BY 0.8 ;
END MAS2796

MACRO MAS2797
   SIZE 1.01 BY 0.8 ;
END MAS2797

MACRO MAS2798
   SIZE 1.01 BY 0.8 ;
END MAS2798

MACRO MAS2799
   SIZE 1.01 BY 0.8 ;
END MAS2799

MACRO MAS2800
   SIZE 1.01 BY 0.8 ;
END MAS2800

MACRO MAS2801
   SIZE 1.01 BY 0.8 ;
END MAS2801

MACRO MAS2802
   SIZE 1.01 BY 0.8 ;
END MAS2802

MACRO MAS2803
   SIZE 1.01 BY 0.8 ;
END MAS2803

MACRO MAS2804
   SIZE 1.01 BY 0.8 ;
END MAS2804

MACRO MAS2805
   SIZE 1.01 BY 0.8 ;
END MAS2805

MACRO MAS2806
   SIZE 1.01 BY 0.8 ;
END MAS2806

MACRO MAS2807
   SIZE 1.01 BY 0.8 ;
END MAS2807

MACRO MAS2808
   SIZE 1.01 BY 0.8 ;
END MAS2808

MACRO MAS2809
   SIZE 1.01 BY 0.8 ;
END MAS2809

MACRO MAS2810
   SIZE 1.01 BY 0.8 ;
END MAS2810

MACRO MAS2811
   SIZE 1.01 BY 0.8 ;
END MAS2811

MACRO MAS2812
   SIZE 1.01 BY 0.8 ;
END MAS2812

MACRO MAS2813
   SIZE 1.01 BY 0.8 ;
END MAS2813

MACRO MAS2814
   SIZE 1.01 BY 0.8 ;
END MAS2814

MACRO MAS2815
   SIZE 1.01 BY 0.8 ;
END MAS2815

MACRO MAS2816
   SIZE 1.01 BY 0.8 ;
END MAS2816

MACRO MAS2817
   SIZE 1.01 BY 0.8 ;
END MAS2817

MACRO MAS2818
   SIZE 1.01 BY 0.8 ;
END MAS2818

MACRO MAS2819
   SIZE 1.01 BY 0.8 ;
END MAS2819

MACRO MAS2820
   SIZE 1.01 BY 0.8 ;
END MAS2820

MACRO MAS2821
   SIZE 1.01 BY 0.8 ;
END MAS2821

MACRO MAS2822
   SIZE 1.01 BY 0.8 ;
END MAS2822

MACRO MAS2823
   SIZE 1.01 BY 0.8 ;
END MAS2823

MACRO MAS2824
   SIZE 1.01 BY 0.8 ;
END MAS2824

MACRO MAS2825
   SIZE 1.01 BY 0.8 ;
END MAS2825

MACRO MAS2826
   SIZE 1.01 BY 0.8 ;
END MAS2826

MACRO MAS2827
   SIZE 1.01 BY 0.8 ;
END MAS2827

MACRO MAS2828
   SIZE 1.01 BY 0.8 ;
END MAS2828

MACRO MAS2829
   SIZE 1.01 BY 0.8 ;
END MAS2829

MACRO MAS2830
   SIZE 1.01 BY 0.8 ;
END MAS2830

MACRO MAS2831
   SIZE 1.01 BY 0.8 ;
END MAS2831

MACRO MAS2832
   SIZE 1.01 BY 0.8 ;
END MAS2832

MACRO MAS2833
   SIZE 1.01 BY 0.8 ;
END MAS2833

MACRO MAS2834
   SIZE 1.01 BY 0.8 ;
END MAS2834

MACRO MAS2835
   SIZE 1.01 BY 0.8 ;
END MAS2835

MACRO MAS2836
   SIZE 1.01 BY 0.8 ;
END MAS2836

MACRO MAS2837
   SIZE 1.01 BY 0.8 ;
END MAS2837

MACRO MAS2838
   SIZE 1.01 BY 0.8 ;
END MAS2838

MACRO MAS2839
   SIZE 1.01 BY 0.8 ;
END MAS2839

MACRO MAS2840
   SIZE 1.01 BY 0.8 ;
END MAS2840

MACRO MAS2841
   SIZE 1.01 BY 0.8 ;
END MAS2841

MACRO MAS2842
   SIZE 1.01 BY 0.8 ;
END MAS2842

MACRO MAS2843
   SIZE 1.1 BY 1.44 ;
END MAS2843

MACRO MAS2844
   SIZE 1.44 BY 1.12 ;
END MAS2844

MACRO MAS2845
   SIZE 7.01 BY 3.84 ;
END MAS2845

