MACRO c0
     SIZE 1056 BY 504 ;
END c0

MACRO c1
     SIZE 924 BY 504 ;
END c1

MACRO c2
     SIZE 792 BY 504 ;
END c2

MACRO c3
     SIZE 132 BY 504 ;
END c3

MACRO c4
     SIZE 396 BY 504 ;
END c4

MACRO c5
     SIZE 528 BY 504 ;
END c5

MACRO c6
     SIZE 264 BY 504 ;
END c6

MACRO c7
     SIZE 1320 BY 504 ;
END c7

MACRO c8
     SIZE 1188 BY 504 ;
END c8

MACRO c9
     SIZE 660 BY 504 ;
END c9

MACRO c10
     SIZE 1584 BY 504 ;
END c10

MACRO c11
     SIZE 1716 BY 504 ;
END c11

MACRO c12
     SIZE 1980 BY 504 ;
END c12

MACRO c13
     SIZE 1848 BY 504 ;
END c13

MACRO c14
     SIZE 1452 BY 504 ;
END c14

MACRO c15
     SIZE 2244 BY 504 ;
END c15

END LIBRARY