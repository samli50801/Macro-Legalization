MACRO block_414x1962_350
   SIZE 157.32 BY 372.78 ;
END block_414x1962_350

MACRO block_341x369_76
   SIZE 129.58 BY 70.11 ;
END block_341x369_76

MACRO block_671x702_95
   SIZE 254.98 BY 133.38 ;
END block_671x702_95

MACRO block_197x171_32
   SIZE 74.86 BY 32.49 ;
END block_197x171_32

MACRO block_189x891_64
   SIZE 71.82 BY 169.29 ;
END block_189x891_64

MACRO block_189x414_32
   SIZE 71.82 BY 78.66 ;
END block_189x414_32

MACRO block_533x5436_977
   SIZE 202.54 BY 1032.84 ;
END block_533x5436_977

MACRO block_416x441_106
   SIZE 158.08 BY 83.79 ;
END block_416x441_106

MACRO block_5572x6435_643
   SIZE 2117.36 BY 1222.65 ;
END block_5572x6435_643

MACRO block_646x2664_73
   SIZE 245.48 BY 506.16 ;
END block_646x2664_73

MACRO block_3700x6435_640
   SIZE 1406.0 BY 1222.65 ;
END block_3700x6435_640

MACRO block_646x2664_74
   SIZE 245.48 BY 506.16 ;
END block_646x2664_74

MACRO block_2456x4212_423
   SIZE 933.28 BY 800.28 ;
END block_2456x4212_423

MACRO block_416x441_112
   SIZE 158.08 BY 83.79 ;
END block_416x441_112

MACRO block_414x2160_386
   SIZE 157.32 BY 410.4 ;
END block_414x2160_386

MACRO block_414x2160_386_1
   SIZE 157.32 BY 410.4 ;
END block_414x2160_386_1

MACRO block_1338x2592_114
   SIZE 508.44 BY 492.48 ;
END block_1338x2592_114

MACRO block_341x369_82
   SIZE 129.58 BY 70.11 ;
END block_341x369_82

MACRO block_779x2592_111
   SIZE 296.02 BY 492.48 ;
END block_779x2592_111

MACRO block_341x369_80
   SIZE 129.58 BY 70.11 ;
END block_341x369_80

MACRO block_535x648_127
   SIZE 203.3 BY 123.12 ;
END block_535x648_127

MACRO block_197x180_32
   SIZE 74.86 BY 34.2 ;
END block_197x180_32

MACRO block_535x648_127_1
   SIZE 203.3 BY 123.12 ;
END block_535x648_127_1

MACRO block_2305x2763_1381
   SIZE 875.9 BY 524.97 ;
END block_2305x2763_1381

MACRO block_336x333_86
   SIZE 127.68 BY 63.27 ;
END block_336x333_86

MACRO block_644x675_97
   SIZE 244.72 BY 128.25 ;
END block_644x675_97

MACRO block_607x549_108
   SIZE 230.66 BY 104.31 ;
END block_607x549_108

MACRO block_607x549_108_1
   SIZE 230.66 BY 104.31 ;
END block_607x549_108_1

MACRO block_535x549_99
   SIZE 203.3 BY 104.31 ;
END block_535x549_99

MACRO block_546x684_108
   SIZE 207.48 BY 129.96 ;
END block_546x684_108

MACRO block_575x315_26
   SIZE 218.5 BY 59.85 ;
END block_575x315_26

MACRO block_96x2439_162
   SIZE 36.48 BY 463.41 ;
END block_96x2439_162

MACRO block_96x1980_132
   SIZE 36.48 BY 376.2 ;
END block_96x1980_132

MACRO block_1338x3105_126
   SIZE 508.44 BY 589.95 ;
END block_1338x3105_126

MACRO block_341x360_82
   SIZE 129.58 BY 68.4 ;
END block_341x360_82

MACRO block_1338x1728_121
   SIZE 508.44 BY 328.32 ;
END block_1338x1728_121

MACRO block_341x369_78
   SIZE 129.58 BY 70.11 ;
END block_341x369_78

MACRO block_535x702_148
   SIZE 203.3 BY 133.38 ;
END block_535x702_148

MACRO block_535x693_148
   SIZE 203.3 BY 131.67 ;
END block_535x693_148

MACRO block_197x180_31
   SIZE 74.86 BY 34.2 ;
END block_197x180_31

MACRO block_2456x2844_180
   SIZE 933.28 BY 540.36 ;
END block_2456x2844_180

MACRO block_341x369_84
   SIZE 129.58 BY 70.11 ;
END block_341x369_84

MACRO block_1338x2844_177
   SIZE 508.44 BY 540.36 ;
END block_1338x2844_177

MACRO block_414x1035_170
   SIZE 157.32 BY 196.65 ;
END block_414x1035_170

MACRO block_341x369_68
   SIZE 129.58 BY 70.11 ;
END block_341x369_68

MACRO block_2456x5499_316
   SIZE 933.28 BY 1044.81 ;
END block_2456x5499_316

MACRO block_546x675_108
   SIZE 207.48 BY 128.25 ;
END block_546x675_108

MACRO block_416x432_112
   SIZE 158.08 BY 82.08 ;
END block_416x432_112

MACRO block_2456x2799_291
   SIZE 933.28 BY 531.81 ;
END block_2456x2799_291

MACRO block_414x1575_274
   SIZE 157.32 BY 299.25 ;
END block_414x1575_274

MACRO block_341x369_72
   SIZE 129.58 BY 70.11 ;
END block_341x369_72

MACRO block_189x648_48
   SIZE 71.82 BY 123.12 ;
END block_189x648_48

MACRO block_414x3861_682
   SIZE 157.32 BY 733.59 ;
END block_414x3861_682

MACRO block_416x441_104
   SIZE 158.08 BY 83.79 ;
END block_416x441_104

MACRO block_546x675_88
   SIZE 207.48 BY 128.25 ;
END block_546x675_88

MACRO block_1338x1728_90
   SIZE 508.44 BY 328.32 ;
END block_1338x1728_90

MACRO block_341x360_78
   SIZE 129.58 BY 68.4 ;
END block_341x360_78

MACRO block_535x549_99_1
   SIZE 203.3 BY 104.31 ;
END block_535x549_99_1

MACRO block_533x1251_217
   SIZE 202.54 BY 237.69 ;
END block_533x1251_217

MACRO block_341x369_74
   SIZE 129.58 BY 70.11 ;
END block_341x369_74

MACRO block_779x2160_225
   SIZE 296.02 BY 410.4 ;
END block_779x2160_225

MACRO block_1829x2160_231
   SIZE 695.02 BY 410.4 ;
END block_1829x2160_231

MACRO block_341x360_84
   SIZE 129.58 BY 68.4 ;
END block_341x360_84

MACRO block_1338x2583_268
   SIZE 508.44 BY 490.77 ;
END block_1338x2583_268

MACRO block_779x1467_260
   SIZE 296.02 BY 278.73 ;
END block_779x1467_260

MACRO block_533x1251_134
   SIZE 202.54 BY 237.69 ;
END block_533x1251_134

MACRO block_1338x1899_98
   SIZE 508.44 BY 360.81 ;
END block_1338x1899_98

MACRO block_546x675_72
   SIZE 207.48 BY 128.25 ;
END block_546x675_72

MACRO block_414x6183_1122
   SIZE 157.32 BY 1174.77 ;
END block_414x6183_1122

MACRO block_779x1107_192
   SIZE 296.02 BY 210.33 ;
END block_779x1107_192

MACRO block_546x675_107
   SIZE 207.48 BY 128.25 ;
END block_546x675_107

MACRO block_341x369_75
   SIZE 129.58 BY 70.11 ;
END block_341x369_75

MACRO block_414x3366_590
   SIZE 157.32 BY 639.54 ;
END block_414x3366_590

MACRO block_414x3438_602
   SIZE 157.32 BY 653.22 ;
END block_414x3438_602

MACRO block_533x1062_181
   SIZE 202.54 BY 201.78 ;
END block_533x1062_181

MACRO block_414x1071_178
   SIZE 157.32 BY 203.49 ;
END block_414x1071_178

MACRO block_126x1134_79
   SIZE 47.88 BY 215.46 ;
END block_126x1134_79

MACRO block_96x1134_78
   SIZE 36.48 BY 215.46 ;
END block_96x1134_78

MACRO block_96x1134_76
   SIZE 36.48 BY 215.46 ;
END block_96x1134_76

MACRO block_533x1062_181_1
   SIZE 202.54 BY 201.78 ;
END block_533x1062_181_1

MACRO block_414x1062_178
   SIZE 157.32 BY 201.78 ;
END block_414x1062_178

MACRO block_126x1134_78
   SIZE 47.88 BY 215.46 ;
END block_126x1134_78

MACRO block_533x1062_181_2
   SIZE 202.54 BY 201.78 ;
END block_533x1062_181_2

MACRO block_546x684_97
   SIZE 207.48 BY 129.96 ;
END block_546x684_97

MACRO block_2456x2763_176
   SIZE 933.28 BY 524.97 ;
END block_2456x2763_176

MACRO block_546x675_92
   SIZE 207.48 BY 128.25 ;
END block_546x675_92

MACRO block_414x1962_350_1
   SIZE 157.32 BY 372.78 ;
END block_414x1962_350_1

MACRO block_341x378_76
   SIZE 129.58 BY 71.82 ;
END block_341x378_76

MACRO block_414x1908_342
   SIZE 157.32 BY 362.52 ;
END block_414x1908_342

MACRO block_341x360_76
   SIZE 129.58 BY 68.4 ;
END block_341x360_76

MACRO block_546x684_98
   SIZE 207.48 BY 129.96 ;
END block_546x684_98

MACRO block_533x1296_225
   SIZE 202.54 BY 246.24 ;
END block_533x1296_225

MACRO block_533x1701_301
   SIZE 202.54 BY 323.19 ;
END block_533x1701_301

MACRO block_341x378_73
   SIZE 129.58 BY 71.82 ;
END block_341x378_73

MACRO block_414x1215_206
   SIZE 157.32 BY 230.85 ;
END block_414x1215_206

MACRO block_535x747_156
   SIZE 203.3 BY 141.93 ;
END block_535x747_156

MACRO block_197x171_33
   SIZE 74.86 BY 32.49 ;
END block_197x171_33

MACRO block_575x315_27
   SIZE 218.5 BY 59.85 ;
END block_575x315_27

MACRO block_779x2223_404
   SIZE 296.02 BY 422.37 ;
END block_779x2223_404

MACRO block_779x1701_304
   SIZE 296.02 BY 323.19 ;
END block_779x1701_304

MACRO block_779x1701_304_1
   SIZE 296.02 BY 323.19 ;
END block_779x1701_304_1

MACRO block_1004x2529_626
   SIZE 381.52 BY 480.51 ;
END block_1004x2529_626

MACRO block_546x675_103
   SIZE 207.48 BY 128.25 ;
END block_546x675_103

MACRO block_232x297_54
   SIZE 88.16 BY 56.43 ;
END block_232x297_54

MACRO block_414x1035_170_1
   SIZE 157.32 BY 196.65 ;
END block_414x1035_170_1

MACRO block_414x3672_646
   SIZE 157.32 BY 697.68 ;
END block_414x3672_646

MACRO block_416x441_103
   SIZE 158.08 BY 83.79 ;
END block_416x441_103

MACRO block_567x648_52
   SIZE 215.46 BY 123.12 ;
END block_567x648_52

MACRO block_567x648_53
   SIZE 215.46 BY 123.12 ;
END block_567x648_53

MACRO block_1829x4383_264
   SIZE 695.02 BY 832.77 ;
END block_1829x4383_264

MACRO block_416x441_111
   SIZE 158.08 BY 83.79 ;
END block_416x441_111

MACRO block_1829x4383_264_1
   SIZE 695.02 BY 832.77 ;
END block_1829x4383_264_1

MACRO block_1829x6012_340
   SIZE 695.02 BY 1142.28 ;
END block_1829x6012_340

MACRO block_546x675_109
   SIZE 207.48 BY 128.25 ;
END block_546x675_109

MACRO block_96x2466_164
   SIZE 36.48 BY 468.54 ;
END block_96x2466_164

MACRO block_323x801_40
   SIZE 122.74 BY 152.19 ;
END block_323x801_40

MACRO block_323x864_42
   SIZE 122.74 BY 164.16 ;
END block_323x864_42

MACRO block_73x72_14
   SIZE 27.74 BY 13.68 ;
END block_73x72_14

MACRO block_73x72_15
   SIZE 27.74 BY 13.68 ;
END block_73x72_15

END LIBRARY
